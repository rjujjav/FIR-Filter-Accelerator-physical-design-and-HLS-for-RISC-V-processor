
//------> /mnt/coe/workspace/ece/ece720-common/tools/catapult2021.1/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /mnt/coe/workspace/ece/ece720-common/tools/catapult2021.1/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> /mnt/coe/workspace/ece/ece720-common/tools/catapult2021.1/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2021.1/950854 Production Release
//  HLS Date:       Mon Aug  2 21:36:02 PDT 2021
// 
//  Generated by:   rjujjav@lib-41917.eos.ncsu.edu
//  Generated date: Sat Dec  9 00:51:56 2023
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Accelerator_run_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module Accelerator_run_run_run_fsm (
  clk, reset_bar, fsm_output, while_C_1_tr0, while_if_for_for_C_0_tr0, while_if_for_C_0_tr0,
      while_if_for_1_for_C_1_tr0, while_if_for_1_C_1_tr0, while_C_2_tr0, while_if_for_2_for_C_1_tr0,
      while_if_for_2_C_1_tr0, while_C_3_tr0, while_if_for_3_for_C_1_tr0, while_if_for_3_C_1_tr0,
      while_C_4_tr0, while_if_for_4_for_C_1_tr0, while_if_for_4_C_1_tr0
);
  input clk;
  input reset_bar;
  output [24:0] fsm_output;
  reg [24:0] fsm_output;
  input while_C_1_tr0;
  input while_if_for_for_C_0_tr0;
  input while_if_for_C_0_tr0;
  input while_if_for_1_for_C_1_tr0;
  input while_if_for_1_C_1_tr0;
  input while_C_2_tr0;
  input while_if_for_2_for_C_1_tr0;
  input while_if_for_2_C_1_tr0;
  input while_C_3_tr0;
  input while_if_for_3_for_C_1_tr0;
  input while_if_for_3_C_1_tr0;
  input while_C_4_tr0;
  input while_if_for_4_for_C_1_tr0;
  input while_if_for_4_C_1_tr0;


  // FSM State Type Declaration for Accelerator_run_run_run_fsm_1
  parameter
    run_rlp_C_0 = 5'd0,
    while_C_0 = 5'd1,
    while_C_1 = 5'd2,
    while_if_for_for_C_0 = 5'd3,
    while_if_for_C_0 = 5'd4,
    while_if_for_1_C_0 = 5'd5,
    while_if_for_1_for_C_0 = 5'd6,
    while_if_for_1_for_C_1 = 5'd7,
    while_if_for_1_C_1 = 5'd8,
    while_C_2 = 5'd9,
    while_if_for_2_C_0 = 5'd10,
    while_if_for_2_for_C_0 = 5'd11,
    while_if_for_2_for_C_1 = 5'd12,
    while_if_for_2_C_1 = 5'd13,
    while_C_3 = 5'd14,
    while_if_for_3_C_0 = 5'd15,
    while_if_for_3_for_C_0 = 5'd16,
    while_if_for_3_for_C_1 = 5'd17,
    while_if_for_3_C_1 = 5'd18,
    while_C_4 = 5'd19,
    while_if_for_4_C_0 = 5'd20,
    while_if_for_4_for_C_0 = 5'd21,
    while_if_for_4_for_C_1 = 5'd22,
    while_if_for_4_C_1 = 5'd23,
    while_C_5 = 5'd24;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : Accelerator_run_run_run_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 25'b0000000000000000000000010;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 25'b0000000000000000000000100;
        if ( while_C_1_tr0 ) begin
          state_var_NS = while_C_2;
        end
        else begin
          state_var_NS = while_if_for_for_C_0;
        end
      end
      while_if_for_for_C_0 : begin
        fsm_output = 25'b0000000000000000000001000;
        if ( while_if_for_for_C_0_tr0 ) begin
          state_var_NS = while_if_for_C_0;
        end
        else begin
          state_var_NS = while_if_for_for_C_0;
        end
      end
      while_if_for_C_0 : begin
        fsm_output = 25'b0000000000000000000010000;
        if ( while_if_for_C_0_tr0 ) begin
          state_var_NS = while_if_for_1_C_0;
        end
        else begin
          state_var_NS = while_if_for_for_C_0;
        end
      end
      while_if_for_1_C_0 : begin
        fsm_output = 25'b0000000000000000000100000;
        state_var_NS = while_if_for_1_for_C_0;
      end
      while_if_for_1_for_C_0 : begin
        fsm_output = 25'b0000000000000000001000000;
        state_var_NS = while_if_for_1_for_C_1;
      end
      while_if_for_1_for_C_1 : begin
        fsm_output = 25'b0000000000000000010000000;
        if ( while_if_for_1_for_C_1_tr0 ) begin
          state_var_NS = while_if_for_1_C_1;
        end
        else begin
          state_var_NS = while_if_for_1_for_C_0;
        end
      end
      while_if_for_1_C_1 : begin
        fsm_output = 25'b0000000000000000100000000;
        if ( while_if_for_1_C_1_tr0 ) begin
          state_var_NS = while_C_2;
        end
        else begin
          state_var_NS = while_if_for_1_C_0;
        end
      end
      while_C_2 : begin
        fsm_output = 25'b0000000000000001000000000;
        if ( while_C_2_tr0 ) begin
          state_var_NS = while_C_3;
        end
        else begin
          state_var_NS = while_if_for_2_C_0;
        end
      end
      while_if_for_2_C_0 : begin
        fsm_output = 25'b0000000000000010000000000;
        state_var_NS = while_if_for_2_for_C_0;
      end
      while_if_for_2_for_C_0 : begin
        fsm_output = 25'b0000000000000100000000000;
        state_var_NS = while_if_for_2_for_C_1;
      end
      while_if_for_2_for_C_1 : begin
        fsm_output = 25'b0000000000001000000000000;
        if ( while_if_for_2_for_C_1_tr0 ) begin
          state_var_NS = while_if_for_2_C_1;
        end
        else begin
          state_var_NS = while_if_for_2_for_C_0;
        end
      end
      while_if_for_2_C_1 : begin
        fsm_output = 25'b0000000000010000000000000;
        if ( while_if_for_2_C_1_tr0 ) begin
          state_var_NS = while_C_3;
        end
        else begin
          state_var_NS = while_if_for_2_C_0;
        end
      end
      while_C_3 : begin
        fsm_output = 25'b0000000000100000000000000;
        if ( while_C_3_tr0 ) begin
          state_var_NS = while_C_4;
        end
        else begin
          state_var_NS = while_if_for_3_C_0;
        end
      end
      while_if_for_3_C_0 : begin
        fsm_output = 25'b0000000001000000000000000;
        state_var_NS = while_if_for_3_for_C_0;
      end
      while_if_for_3_for_C_0 : begin
        fsm_output = 25'b0000000010000000000000000;
        state_var_NS = while_if_for_3_for_C_1;
      end
      while_if_for_3_for_C_1 : begin
        fsm_output = 25'b0000000100000000000000000;
        if ( while_if_for_3_for_C_1_tr0 ) begin
          state_var_NS = while_if_for_3_C_1;
        end
        else begin
          state_var_NS = while_if_for_3_for_C_0;
        end
      end
      while_if_for_3_C_1 : begin
        fsm_output = 25'b0000001000000000000000000;
        if ( while_if_for_3_C_1_tr0 ) begin
          state_var_NS = while_C_4;
        end
        else begin
          state_var_NS = while_if_for_3_C_0;
        end
      end
      while_C_4 : begin
        fsm_output = 25'b0000010000000000000000000;
        if ( while_C_4_tr0 ) begin
          state_var_NS = while_C_5;
        end
        else begin
          state_var_NS = while_if_for_4_C_0;
        end
      end
      while_if_for_4_C_0 : begin
        fsm_output = 25'b0000100000000000000000000;
        state_var_NS = while_if_for_4_for_C_0;
      end
      while_if_for_4_for_C_0 : begin
        fsm_output = 25'b0001000000000000000000000;
        state_var_NS = while_if_for_4_for_C_1;
      end
      while_if_for_4_for_C_1 : begin
        fsm_output = 25'b0010000000000000000000000;
        if ( while_if_for_4_for_C_1_tr0 ) begin
          state_var_NS = while_if_for_4_C_1;
        end
        else begin
          state_var_NS = while_if_for_4_for_C_0;
        end
      end
      while_if_for_4_C_1 : begin
        fsm_output = 25'b0100000000000000000000000;
        if ( while_if_for_4_C_1_tr0 ) begin
          state_var_NS = while_C_5;
        end
        else begin
          state_var_NS = while_if_for_4_C_0;
        end
      end
      while_C_5 : begin
        fsm_output = 25'b1000000000000000000000000;
        state_var_NS = while_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 25'b0000000000000000000000001;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      state_var <= run_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_run_fsm (
  clk, reset_bar, run_wen, fsm_output
);
  input clk;
  input reset_bar;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for AxiSlaveToReg2_axi_cfg_standard_14_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : AxiSlaveToReg2_axi_cfg_standard_14_16_run_run_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_staller
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_staller (
  clk, reset_bar, run_wen, run_wten, if_axi_rd_r_Push_mioi_wen_comp, if_axi_wr_b_Push_mioi_wen_comp,
      run_flen_unreg
);
  input clk;
  input reset_bar;
  output run_wen;
  output run_wten;
  reg run_wten;
  input if_axi_rd_r_Push_mioi_wen_comp;
  input if_axi_wr_b_Push_mioi_wen_comp;
  input run_flen_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = if_axi_rd_r_Push_mioi_wen_comp & if_axi_wr_b_Push_mioi_wen_comp
      & (~ run_flen_unreg);
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      run_wten <= 1'b0;
    end
    else begin
      run_wten <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_if_axi_wr_b_Push_mio_wait_dp
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_if_axi_wr_b_Push_mio_wait_dp
    (
  clk, reset_bar, if_axi_wr_b_Push_mioi_oswt_unreg, if_axi_wr_b_Push_mioi_bawt, if_axi_wr_b_Push_mioi_wen_comp,
      if_axi_wr_b_Push_mioi_biwt, if_axi_wr_b_Push_mioi_bdwt
);
  input clk;
  input reset_bar;
  input if_axi_wr_b_Push_mioi_oswt_unreg;
  output if_axi_wr_b_Push_mioi_bawt;
  output if_axi_wr_b_Push_mioi_wen_comp;
  input if_axi_wr_b_Push_mioi_biwt;
  input if_axi_wr_b_Push_mioi_bdwt;


  // Interconnect Declarations
  reg if_axi_wr_b_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign if_axi_wr_b_Push_mioi_bawt = if_axi_wr_b_Push_mioi_biwt | if_axi_wr_b_Push_mioi_bcwt;
  assign if_axi_wr_b_Push_mioi_wen_comp = (~ if_axi_wr_b_Push_mioi_oswt_unreg) |
      if_axi_wr_b_Push_mioi_bawt;
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_b_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      if_axi_wr_b_Push_mioi_bcwt <= ~((~(if_axi_wr_b_Push_mioi_bcwt | if_axi_wr_b_Push_mioi_biwt))
          | if_axi_wr_b_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_if_axi_wr_b_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_if_axi_wr_b_Push_mio_wait_ctrl
    (
  clk, reset_bar, run_wen, run_wten, if_axi_wr_b_Push_mioi_oswt_unreg, if_axi_wr_b_Push_mioi_iswt0,
      if_axi_wr_b_Push_mioi_biwt, if_axi_wr_b_Push_mioi_bdwt, if_axi_wr_b_Push_mioi_ivld_run_sct,
      if_axi_wr_b_Push_mioi_irdy
);
  input clk;
  input reset_bar;
  input run_wen;
  input run_wten;
  input if_axi_wr_b_Push_mioi_oswt_unreg;
  input if_axi_wr_b_Push_mioi_iswt0;
  output if_axi_wr_b_Push_mioi_biwt;
  output if_axi_wr_b_Push_mioi_bdwt;
  output if_axi_wr_b_Push_mioi_ivld_run_sct;
  input if_axi_wr_b_Push_mioi_irdy;


  // Interconnect Declarations
  wire if_axi_wr_b_Push_mioi_ogwt;
  reg if_axi_wr_b_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign if_axi_wr_b_Push_mioi_bdwt = if_axi_wr_b_Push_mioi_oswt_unreg & run_wen;
  assign if_axi_wr_b_Push_mioi_biwt = if_axi_wr_b_Push_mioi_ogwt & if_axi_wr_b_Push_mioi_irdy;
  assign if_axi_wr_b_Push_mioi_ogwt = ((~ run_wten) & if_axi_wr_b_Push_mioi_iswt0)
      | if_axi_wr_b_Push_mioi_icwt;
  assign if_axi_wr_b_Push_mioi_ivld_run_sct = if_axi_wr_b_Push_mioi_ogwt;
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_b_Push_mioi_icwt <= 1'b0;
    end
    else begin
      if_axi_wr_b_Push_mioi_icwt <= if_axi_wr_b_Push_mioi_ogwt & (~ if_axi_wr_b_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_if_axi_wr_w_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_if_axi_wr_w_PopNB_mio_wait_dp
    (
  clk, reset_bar, if_axi_wr_w_PopNB_mioi_bawt, if_axi_wr_w_PopNB_mioi_ivld_mxwt,
      if_axi_wr_w_PopNB_mioi_idat_mxwt, if_axi_wr_w_PopNB_mioi_biwt, if_axi_wr_w_PopNB_mioi_bdwt,
      if_axi_wr_w_PopNB_mioi_ivld, if_axi_wr_w_PopNB_mioi_idat
);
  input clk;
  input reset_bar;
  output if_axi_wr_w_PopNB_mioi_bawt;
  output if_axi_wr_w_PopNB_mioi_ivld_mxwt;
  output [72:0] if_axi_wr_w_PopNB_mioi_idat_mxwt;
  input if_axi_wr_w_PopNB_mioi_biwt;
  input if_axi_wr_w_PopNB_mioi_bdwt;
  input if_axi_wr_w_PopNB_mioi_ivld;
  input [72:0] if_axi_wr_w_PopNB_mioi_idat;


  // Interconnect Declarations
  reg if_axi_wr_w_PopNB_mioi_bcwt;
  reg if_axi_wr_w_PopNB_mioi_ivld_bfwt;
  reg [72:0] if_axi_wr_w_PopNB_mioi_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign if_axi_wr_w_PopNB_mioi_bawt = if_axi_wr_w_PopNB_mioi_biwt | if_axi_wr_w_PopNB_mioi_bcwt;
  assign if_axi_wr_w_PopNB_mioi_ivld_mxwt = MUX_s_1_2_2(if_axi_wr_w_PopNB_mioi_ivld,
      if_axi_wr_w_PopNB_mioi_ivld_bfwt, if_axi_wr_w_PopNB_mioi_bcwt);
  assign if_axi_wr_w_PopNB_mioi_idat_mxwt = MUX_v_73_2_2(if_axi_wr_w_PopNB_mioi_idat,
      if_axi_wr_w_PopNB_mioi_idat_bfwt, if_axi_wr_w_PopNB_mioi_bcwt);
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_w_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      if_axi_wr_w_PopNB_mioi_bcwt <= ~((~(if_axi_wr_w_PopNB_mioi_bcwt | if_axi_wr_w_PopNB_mioi_biwt))
          | if_axi_wr_w_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_w_PopNB_mioi_ivld_bfwt <= 1'b0;
      if_axi_wr_w_PopNB_mioi_idat_bfwt <= 73'b0000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( if_axi_wr_w_PopNB_mioi_biwt ) begin
      if_axi_wr_w_PopNB_mioi_ivld_bfwt <= if_axi_wr_w_PopNB_mioi_ivld;
      if_axi_wr_w_PopNB_mioi_idat_bfwt <= if_axi_wr_w_PopNB_mioi_idat;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [72:0] MUX_v_73_2_2;
    input [72:0] input_0;
    input [72:0] input_1;
    input  sel;
    reg [72:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_73_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_if_axi_wr_w_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_if_axi_wr_w_PopNB_mio_wait_ctrl
    (
  run_wen, run_wten, if_axi_wr_w_PopNB_mioi_oswt_unreg, if_axi_wr_w_PopNB_mioi_iswt0,
      if_axi_wr_w_PopNB_mioi_biwt, if_axi_wr_w_PopNB_mioi_bdwt
);
  input run_wen;
  input run_wten;
  input if_axi_wr_w_PopNB_mioi_oswt_unreg;
  input if_axi_wr_w_PopNB_mioi_iswt0;
  output if_axi_wr_w_PopNB_mioi_biwt;
  output if_axi_wr_w_PopNB_mioi_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign if_axi_wr_w_PopNB_mioi_bdwt = if_axi_wr_w_PopNB_mioi_oswt_unreg & run_wen;
  assign if_axi_wr_w_PopNB_mioi_biwt = (~ run_wten) & if_axi_wr_w_PopNB_mioi_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_if_axi_rd_r_Push_mio_wait_dp
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_if_axi_rd_r_Push_mio_wait_dp
    (
  clk, reset_bar, if_axi_rd_r_Push_mioi_oswt_unreg, if_axi_rd_r_Push_mioi_bawt, if_axi_rd_r_Push_mioi_wen_comp,
      if_axi_rd_r_Push_mioi_biwt, if_axi_rd_r_Push_mioi_bdwt
);
  input clk;
  input reset_bar;
  input if_axi_rd_r_Push_mioi_oswt_unreg;
  output if_axi_rd_r_Push_mioi_bawt;
  output if_axi_rd_r_Push_mioi_wen_comp;
  input if_axi_rd_r_Push_mioi_biwt;
  input if_axi_rd_r_Push_mioi_bdwt;


  // Interconnect Declarations
  reg if_axi_rd_r_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign if_axi_rd_r_Push_mioi_bawt = if_axi_rd_r_Push_mioi_biwt | if_axi_rd_r_Push_mioi_bcwt;
  assign if_axi_rd_r_Push_mioi_wen_comp = (~ if_axi_rd_r_Push_mioi_oswt_unreg) |
      if_axi_rd_r_Push_mioi_bawt;
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_rd_r_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      if_axi_rd_r_Push_mioi_bcwt <= ~((~(if_axi_rd_r_Push_mioi_bcwt | if_axi_rd_r_Push_mioi_biwt))
          | if_axi_rd_r_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_if_axi_rd_r_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_if_axi_rd_r_Push_mio_wait_ctrl
    (
  clk, reset_bar, run_wen, run_wten, if_axi_rd_r_Push_mioi_oswt_unreg, if_axi_rd_r_Push_mioi_iswt0,
      if_axi_rd_r_Push_mioi_biwt, if_axi_rd_r_Push_mioi_bdwt, if_axi_rd_r_Push_mioi_ivld_run_sct,
      if_axi_rd_r_Push_mioi_irdy
);
  input clk;
  input reset_bar;
  input run_wen;
  input run_wten;
  input if_axi_rd_r_Push_mioi_oswt_unreg;
  input if_axi_rd_r_Push_mioi_iswt0;
  output if_axi_rd_r_Push_mioi_biwt;
  output if_axi_rd_r_Push_mioi_bdwt;
  output if_axi_rd_r_Push_mioi_ivld_run_sct;
  input if_axi_rd_r_Push_mioi_irdy;


  // Interconnect Declarations
  wire if_axi_rd_r_Push_mioi_ogwt;
  reg if_axi_rd_r_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign if_axi_rd_r_Push_mioi_bdwt = if_axi_rd_r_Push_mioi_oswt_unreg & run_wen;
  assign if_axi_rd_r_Push_mioi_biwt = if_axi_rd_r_Push_mioi_ogwt & if_axi_rd_r_Push_mioi_irdy;
  assign if_axi_rd_r_Push_mioi_ogwt = ((~ run_wten) & if_axi_rd_r_Push_mioi_iswt0)
      | if_axi_rd_r_Push_mioi_icwt;
  assign if_axi_rd_r_Push_mioi_ivld_run_sct = if_axi_rd_r_Push_mioi_ogwt;
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_rd_r_Push_mioi_icwt <= 1'b0;
    end
    else begin
      if_axi_rd_r_Push_mioi_icwt <= if_axi_rd_r_Push_mioi_ogwt & (~ if_axi_rd_r_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_regIn_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_regIn_PopNB_mio_wait_dp
    (
  clk, reset_bar, regIn_PopNB_mioi_bawt, regIn_PopNB_mioi_ivld_mxwt, regIn_PopNB_mioi_idat_mxwt,
      regIn_PopNB_mioi_biwt, regIn_PopNB_mioi_bdwt, regIn_PopNB_mioi_ivld, regIn_PopNB_mioi_idat
);
  input clk;
  input reset_bar;
  output regIn_PopNB_mioi_bawt;
  output regIn_PopNB_mioi_ivld_mxwt;
  output [67:0] regIn_PopNB_mioi_idat_mxwt;
  input regIn_PopNB_mioi_biwt;
  input regIn_PopNB_mioi_bdwt;
  input regIn_PopNB_mioi_ivld;
  input [70:0] regIn_PopNB_mioi_idat;


  // Interconnect Declarations
  reg regIn_PopNB_mioi_bcwt;
  reg regIn_PopNB_mioi_ivld_bfwt;
  reg [67:0] regIn_PopNB_mioi_idat_bfwt_70_3;


  // Interconnect Declarations for Component Instantiations 
  assign regIn_PopNB_mioi_bawt = regIn_PopNB_mioi_biwt | regIn_PopNB_mioi_bcwt;
  assign regIn_PopNB_mioi_ivld_mxwt = MUX_s_1_2_2(regIn_PopNB_mioi_ivld, regIn_PopNB_mioi_ivld_bfwt,
      regIn_PopNB_mioi_bcwt);
  assign regIn_PopNB_mioi_idat_mxwt = MUX_v_68_2_2((regIn_PopNB_mioi_idat[70:3]),
      regIn_PopNB_mioi_idat_bfwt_70_3, regIn_PopNB_mioi_bcwt);
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regIn_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      regIn_PopNB_mioi_bcwt <= ~((~(regIn_PopNB_mioi_bcwt | regIn_PopNB_mioi_biwt))
          | regIn_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regIn_PopNB_mioi_ivld_bfwt <= 1'b0;
      regIn_PopNB_mioi_idat_bfwt_70_3 <= 68'b00000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( regIn_PopNB_mioi_biwt ) begin
      regIn_PopNB_mioi_ivld_bfwt <= regIn_PopNB_mioi_ivld;
      regIn_PopNB_mioi_idat_bfwt_70_3 <= regIn_PopNB_mioi_idat[70:3];
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [67:0] MUX_v_68_2_2;
    input [67:0] input_0;
    input [67:0] input_1;
    input  sel;
    reg [67:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_68_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_regIn_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_regIn_PopNB_mio_wait_ctrl
    (
  run_wen, run_wten, regIn_PopNB_mioi_oswt_unreg, regIn_PopNB_mioi_iswt0, regIn_PopNB_mioi_biwt,
      regIn_PopNB_mioi_bdwt
);
  input run_wen;
  input run_wten;
  input regIn_PopNB_mioi_oswt_unreg;
  input regIn_PopNB_mioi_iswt0;
  output regIn_PopNB_mioi_biwt;
  output regIn_PopNB_mioi_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign regIn_PopNB_mioi_bdwt = regIn_PopNB_mioi_oswt_unreg & run_wen;
  assign regIn_PopNB_mioi_biwt = (~ run_wten) & regIn_PopNB_mioi_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_if_axi_wr_aw_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_if_axi_wr_aw_PopNB_mio_wait_dp
    (
  clk, reset_bar, if_axi_wr_aw_PopNB_mioi_bawt, if_axi_wr_aw_PopNB_mioi_ivld_mxwt,
      if_axi_wr_aw_PopNB_mioi_idat_mxwt, if_axi_wr_aw_PopNB_mioi_biwt, if_axi_wr_aw_PopNB_mioi_bdwt,
      if_axi_wr_aw_PopNB_mioi_ivld, if_axi_wr_aw_PopNB_mioi_idat
);
  input clk;
  input reset_bar;
  output if_axi_wr_aw_PopNB_mioi_bawt;
  output if_axi_wr_aw_PopNB_mioi_ivld_mxwt;
  output [19:0] if_axi_wr_aw_PopNB_mioi_idat_mxwt;
  input if_axi_wr_aw_PopNB_mioi_biwt;
  input if_axi_wr_aw_PopNB_mioi_bdwt;
  input if_axi_wr_aw_PopNB_mioi_ivld;
  input [43:0] if_axi_wr_aw_PopNB_mioi_idat;


  // Interconnect Declarations
  reg if_axi_wr_aw_PopNB_mioi_bcwt;
  reg if_axi_wr_aw_PopNB_mioi_ivld_bfwt;
  reg [19:0] if_axi_wr_aw_PopNB_mioi_idat_bfwt_19_0;


  // Interconnect Declarations for Component Instantiations 
  assign if_axi_wr_aw_PopNB_mioi_bawt = if_axi_wr_aw_PopNB_mioi_biwt | if_axi_wr_aw_PopNB_mioi_bcwt;
  assign if_axi_wr_aw_PopNB_mioi_ivld_mxwt = MUX_s_1_2_2(if_axi_wr_aw_PopNB_mioi_ivld,
      if_axi_wr_aw_PopNB_mioi_ivld_bfwt, if_axi_wr_aw_PopNB_mioi_bcwt);
  assign if_axi_wr_aw_PopNB_mioi_idat_mxwt = MUX_v_20_2_2((if_axi_wr_aw_PopNB_mioi_idat[19:0]),
      if_axi_wr_aw_PopNB_mioi_idat_bfwt_19_0, if_axi_wr_aw_PopNB_mioi_bcwt);
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_aw_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      if_axi_wr_aw_PopNB_mioi_bcwt <= ~((~(if_axi_wr_aw_PopNB_mioi_bcwt | if_axi_wr_aw_PopNB_mioi_biwt))
          | if_axi_wr_aw_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_aw_PopNB_mioi_ivld_bfwt <= 1'b0;
      if_axi_wr_aw_PopNB_mioi_idat_bfwt_19_0 <= 20'b00000000000000000000;
    end
    else if ( if_axi_wr_aw_PopNB_mioi_biwt ) begin
      if_axi_wr_aw_PopNB_mioi_ivld_bfwt <= if_axi_wr_aw_PopNB_mioi_ivld;
      if_axi_wr_aw_PopNB_mioi_idat_bfwt_19_0 <= if_axi_wr_aw_PopNB_mioi_idat[19:0];
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_if_axi_wr_aw_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_if_axi_wr_aw_PopNB_mio_wait_ctrl
    (
  run_wen, run_wten, if_axi_wr_aw_PopNB_mioi_oswt_unreg, if_axi_wr_aw_PopNB_mioi_iswt0,
      if_axi_wr_aw_PopNB_mioi_biwt, if_axi_wr_aw_PopNB_mioi_bdwt
);
  input run_wen;
  input run_wten;
  input if_axi_wr_aw_PopNB_mioi_oswt_unreg;
  input if_axi_wr_aw_PopNB_mioi_iswt0;
  output if_axi_wr_aw_PopNB_mioi_biwt;
  output if_axi_wr_aw_PopNB_mioi_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign if_axi_wr_aw_PopNB_mioi_bdwt = if_axi_wr_aw_PopNB_mioi_oswt_unreg & run_wen;
  assign if_axi_wr_aw_PopNB_mioi_biwt = (~ run_wten) & if_axi_wr_aw_PopNB_mioi_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_if_axi_rd_ar_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_if_axi_rd_ar_PopNB_mio_wait_dp
    (
  clk, reset_bar, if_axi_rd_ar_PopNB_mioi_bawt, if_axi_rd_ar_PopNB_mioi_ivld_mxwt,
      if_axi_rd_ar_PopNB_mioi_idat_mxwt, if_axi_rd_ar_PopNB_mioi_biwt, if_axi_rd_ar_PopNB_mioi_bdwt,
      if_axi_rd_ar_PopNB_mioi_ivld, if_axi_rd_ar_PopNB_mioi_idat
);
  input clk;
  input reset_bar;
  output if_axi_rd_ar_PopNB_mioi_bawt;
  output if_axi_rd_ar_PopNB_mioi_ivld_mxwt;
  output [27:0] if_axi_rd_ar_PopNB_mioi_idat_mxwt;
  input if_axi_rd_ar_PopNB_mioi_biwt;
  input if_axi_rd_ar_PopNB_mioi_bdwt;
  input if_axi_rd_ar_PopNB_mioi_ivld;
  input [43:0] if_axi_rd_ar_PopNB_mioi_idat;


  // Interconnect Declarations
  reg if_axi_rd_ar_PopNB_mioi_bcwt;
  reg if_axi_rd_ar_PopNB_mioi_ivld_bfwt;
  reg [43:0] if_axi_rd_ar_PopNB_mioi_idat_bfwt;
  wire [43:0] if_axi_rd_ar_PopNB_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  assign if_axi_rd_ar_PopNB_mioi_bawt = if_axi_rd_ar_PopNB_mioi_biwt | if_axi_rd_ar_PopNB_mioi_bcwt;
  assign if_axi_rd_ar_PopNB_mioi_ivld_mxwt = MUX_s_1_2_2(if_axi_rd_ar_PopNB_mioi_ivld,
      if_axi_rd_ar_PopNB_mioi_ivld_bfwt, if_axi_rd_ar_PopNB_mioi_bcwt);
  assign if_axi_rd_ar_PopNB_mioi_idat_mxwt_pconst = MUX_v_44_2_2(if_axi_rd_ar_PopNB_mioi_idat,
      if_axi_rd_ar_PopNB_mioi_idat_bfwt, if_axi_rd_ar_PopNB_mioi_bcwt);
  assign if_axi_rd_ar_PopNB_mioi_idat_mxwt = {(if_axi_rd_ar_PopNB_mioi_idat_mxwt_pconst[43:36])
      , (if_axi_rd_ar_PopNB_mioi_idat_mxwt_pconst[19:0])};
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_rd_ar_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      if_axi_rd_ar_PopNB_mioi_bcwt <= ~((~(if_axi_rd_ar_PopNB_mioi_bcwt | if_axi_rd_ar_PopNB_mioi_biwt))
          | if_axi_rd_ar_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_rd_ar_PopNB_mioi_ivld_bfwt <= 1'b0;
      if_axi_rd_ar_PopNB_mioi_idat_bfwt <= 44'b00000000000000000000000000000000000000000000;
    end
    else if ( if_axi_rd_ar_PopNB_mioi_biwt ) begin
      if_axi_rd_ar_PopNB_mioi_ivld_bfwt <= if_axi_rd_ar_PopNB_mioi_ivld;
      if_axi_rd_ar_PopNB_mioi_idat_bfwt <= if_axi_rd_ar_PopNB_mioi_idat;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [43:0] MUX_v_44_2_2;
    input [43:0] input_0;
    input [43:0] input_1;
    input  sel;
    reg [43:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_44_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_if_axi_rd_ar_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_if_axi_rd_ar_PopNB_mio_wait_ctrl
    (
  run_wen, run_wten, if_axi_rd_ar_PopNB_mioi_oswt_unreg, if_axi_rd_ar_PopNB_mioi_iswt0,
      if_axi_rd_ar_PopNB_mioi_biwt, if_axi_rd_ar_PopNB_mioi_bdwt
);
  input run_wen;
  input run_wten;
  input if_axi_rd_ar_PopNB_mioi_oswt_unreg;
  input if_axi_rd_ar_PopNB_mioi_iswt0;
  output if_axi_rd_ar_PopNB_mioi_biwt;
  output if_axi_rd_ar_PopNB_mioi_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign if_axi_rd_ar_PopNB_mioi_bdwt = if_axi_rd_ar_PopNB_mioi_oswt_unreg & run_wen;
  assign if_axi_rd_ar_PopNB_mioi_biwt = (~ run_wten) & if_axi_rd_ar_PopNB_mioi_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Accelerator_run_run
// ------------------------------------------------------------------


module Accelerator_run_run (
  clk, reset_bar, regOut_chan_1, regOut_chan_2, regOut_chan_3, regOut_chan_4, regOut_chan_5,
      regOut_chan_6, regOut_chan_7, regOut_chan_8, regOut_chan_9, regIn_chan_PushNB_mioi_ivld,
      regIn_chan_PushNB_mioi_irdy, regIn_chan_PushNB_mioi_idat
);
  input clk;
  input reset_bar;
  input [63:0] regOut_chan_1;
  input [63:0] regOut_chan_2;
  input [63:0] regOut_chan_3;
  input [63:0] regOut_chan_4;
  input [63:0] regOut_chan_5;
  input [63:0] regOut_chan_6;
  input [63:0] regOut_chan_7;
  input [63:0] regOut_chan_8;
  input [63:0] regOut_chan_9;
  output regIn_chan_PushNB_mioi_ivld;
  reg regIn_chan_PushNB_mioi_ivld;
  input regIn_chan_PushNB_mioi_irdy;
  output [70:0] regIn_chan_PushNB_mioi_idat;


  // Interconnect Declarations
  wire [24:0] fsm_output;
  wire [3:0] while_if_for_2_for_1_acc_1_tmp;
  wire [4:0] nl_while_if_for_2_for_1_acc_1_tmp;
  wire while_if_nor_1_tmp;
  wire operator_64_false_1_nor_tmp;
  wire and_dcpl_1;
  wire and_dcpl_3;
  wire or_dcpl_55;
  wire and_dcpl_37;
  wire or_dcpl_135;
  wire or_dcpl_136;
  wire or_dcpl_139;
  wire or_dcpl_142;
  wire or_dcpl_144;
  wire or_dcpl_150;
  wire and_dcpl_55;
  wire and_dcpl_58;
  wire or_dcpl_165;
  wire and_dcpl_61;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_69;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire and_dcpl_78;
  wire or_dcpl_204;
  wire or_dcpl_208;
  wire or_dcpl_209;
  wire or_tmp_141;
  wire or_tmp_197;
  wire or_tmp_331;
  wire or_tmp_333;
  wire and_189_cse;
  wire and_219_cse;
  wire and_225_cse;
  wire and_707_cse;
  wire and_842_cse;
  reg exit_while_if_for_1_for_1_sva;
  reg while_lor_lpi_1_dfm_st;
  reg while_if_for_4_and_tmp_2_sva;
  reg [2:0] while_if_for_4_acc_1_cse_1_sva;
  reg [1:0] while_if_for_1_j_2_0_sva_1_0;
  reg while_if_for_4_and_tmp_1_sva;
  reg while_if_for_4_and_tmp_sva;
  reg [1:0] while_if_for_for_b_2_0_sva_1_0;
  reg [3:0] while_if_for_1_for_1_n_3_0_sva;
  wire regIn_chan_fifo_write_push_mux_1_cse;
  wire regIn_chan_fifo_write_incrHead_mux_cse;
  wire regIn_chan_fifo_write_push_1_mux_1_cse;
  wire regIn_chan_fifo_write_incrHead_1_mux_cse;
  wire regIn_chan_fifo_write_push_2_mux_1_cse;
  wire regIn_chan_fifo_write_incrHead_2_mux_cse;
  wire regIn_chan_fifo_write_push_3_mux_1_cse;
  wire regIn_chan_fifo_write_incrHead_3_mux_cse;
  wire regIn_chan_fifo_write_push_4_mux_1_cse;
  wire regIn_chan_fifo_write_incrHead_4_mux_cse;
  wire or_165_cse;
  wire [15:0] while_if_for_1_and_5_cse;
  wire nand_11_cse;
  wire [15:0] while_if_for_1_and_4_cse;
  wire mux_1_cse;
  wire while_if_for_1_while_if_for_1_or_1_cse;
  reg [63:0] reg_regIn_chan_PushNB_mioi_idat_ftd;
  wire in_equal_cse;
  wire in_equal_1_cse;
  wire in_equal_2_cse;
  wire in_equal_3_cse;
  wire and_107_cse;
  reg [15:0] out_0_lpi_2;
  reg [15:0] out_1_lpi_2;
  reg [15:0] while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva;
  wire [16:0] nl_while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva;
  reg [15:0] out_12_sva;
  wire [4:0] z_out;
  wire [5:0] nl_z_out;
  wire [63:0] z_out_3;
  wire [15:0] z_out_4;
  reg [15:0] we_7_sva;
  reg [15:0] we_8_sva;
  reg [15:0] we_6_sva;
  reg [15:0] we_9_sva;
  reg [15:0] we_5_sva;
  reg [15:0] we_10_sva;
  reg [15:0] we_4_sva;
  reg [15:0] we_11_sva;
  reg [15:0] we_3_sva;
  reg [15:0] we_12_sva;
  reg [15:0] we_2_sva;
  reg [15:0] we_13_sva;
  reg [15:0] we_1_sva;
  reg [15:0] we_14_sva;
  reg [15:0] we_15_sva;
  reg [15:0] in_7_sva;
  reg [15:0] in_8_sva;
  reg [15:0] in_6_sva;
  reg [15:0] in_9_sva;
  reg [15:0] in_5_sva;
  reg [15:0] in_10_sva;
  reg [15:0] in_4_sva;
  reg [15:0] in_11_sva;
  reg [15:0] in_3_sva;
  reg [15:0] in_12_sva;
  reg [15:0] in_2_sva;
  reg [15:0] in_13_sva;
  reg [15:0] in_1_sva;
  reg [15:0] in_14_sva;
  reg [15:0] in_0_sva;
  reg [15:0] out_7_sva;
  reg [15:0] out_6_sva;
  reg [15:0] out_9_sva;
  reg [15:0] out_5_sva;
  reg [15:0] out_10_sva;
  reg [15:0] out_11_sva;
  reg [15:0] out_3_sva;
  reg [15:0] out_2_sva;
  reg [15:0] out_1_sva;
  reg regIn_chan_fifo_write_valid_1_sva;
  reg [15:0] out_10_lpi_2;
  reg [15:0] out_11_lpi_2;
  reg [15:0] we_7_lpi_3;
  reg [15:0] we_8_lpi_3;
  reg [15:0] we_6_lpi_3;
  reg [15:0] we_9_lpi_3;
  reg [15:0] we_5_lpi_3;
  reg [15:0] we_10_lpi_3;
  reg [15:0] we_4_lpi_3;
  reg [15:0] we_11_lpi_3;
  reg [15:0] we_3_lpi_3;
  reg [15:0] we_12_lpi_3;
  reg [15:0] we_2_lpi_3;
  reg [15:0] we_13_lpi_3;
  reg [15:0] we_1_lpi_3;
  reg [15:0] we_14_lpi_3;
  reg [15:0] we_0_lpi_3;
  reg [15:0] we_15_lpi_3;
  reg [63:0] regwr_data_1_sva;
  reg [15:0] in_7_lpi_3;
  reg [15:0] in_8_lpi_3;
  reg [15:0] in_6_lpi_3;
  reg [15:0] in_9_lpi_3;
  reg [15:0] in_5_lpi_3;
  reg [15:0] in_10_lpi_3;
  reg [15:0] in_4_lpi_3;
  reg [15:0] in_11_lpi_3;
  reg [15:0] in_3_lpi_3;
  reg [15:0] in_12_lpi_3;
  reg [15:0] in_2_lpi_3;
  reg [15:0] in_13_lpi_3;
  reg [15:0] in_1_lpi_3;
  reg [15:0] in_14_lpi_3;
  reg [15:0] in_0_lpi_3;
  reg [15:0] in_15_1_sva;
  reg [15:0] out_3_sva_1;
  reg [15:0] out_2_sva_1;
  reg [15:0] out_1_sva_1;
  reg regIn_chan_TransferNBWrite_1_if_asn_mdf_sva;
  reg [15:0] out_7_sva_1;
  reg [15:0] out_6_sva_1;
  reg [15:0] out_5_sva_1;
  wire [15:0] out_3_sva_1_mx0w0;
  wire [15:0] operator_64_false_rshift_ctmp_sva_2;
  wire operator_64_false_nor_m1c_1;
  wire operator_64_false_and_m1c_3;
  wire operator_64_false_and_m1c_4;
  wire operator_64_false_and_m1c_5;
  wire regwr_data_1_sva_mx0c0;
  wire [63:0] regwr_data_1_sva_2;
  wire [15:0] while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1;
  wire while_if_for_4_and_tmp_sva_mx0w0;
  wire while_if_for_4_and_tmp_1_sva_mx0w0;
  wire while_if_for_4_and_tmp_2_sva_mx0w0;
  wire [15:0] while_if_for_1_for_mux_38;
  wire [15:0] while_if_for_2_for_while_if_for_2_for_mux_2;
  wire [15:0] while_if_for_1_for_mul_2;
  wire signed [31:0] nl_while_if_for_1_for_mul_2;
  wire or_601_ssc;
  wire out_or_cse;
  wire and_tmp;
  wire or_tmp_432;
  wire or_tmp_433;
  wire mux_tmp_36;
  wire [4:0] while_if_for_1_for_m_mux_1_rgt;
  reg while_if_for_1_for_m_4_0_sva_1_4;
  reg [3:0] while_if_for_1_for_m_4_0_sva_1_3_0;
  wire and_919_cse;
  wire and_508_cse;
  wire or_636_cse;
  wire or_633_cse;
  wire nand_19_cse;
  wire or_629_cse;
  wire and_753_cse;
  wire and_774_cse;
  wire or_716_cse;
  wire nor_104_cse;
  wire and_809_cse;
  wire or_619_cse;
  reg reg_regIn_chan_PushNB_mioi_idat_1_ftd_3;
  reg [2:0] reg_regIn_chan_PushNB_mioi_idat_1_ftd_2_0;

  wire p_isFull_Pushing_data_to_full_FIFO_prb;
  wire p_isFull_Pushing_data_to_full_FIFO_ctrl_prb;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_prb;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb;
  wire and_104_nl;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_prb;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb;
  wire p_isFull_Pushing_data_to_full_FIFO_prb_1;
  wire p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_1;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_prb_1;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_1;
  wire and_217_nl;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_prb_1;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_1;
  wire p_isFull_Pushing_data_to_full_FIFO_prb_2;
  wire p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_2;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_prb_2;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_2;
  wire and_223_nl;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_prb_2;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_2;
  wire p_isFull_Pushing_data_to_full_FIFO_prb_3;
  wire p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_3;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_prb_3;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_3;
  wire and_229_nl;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_prb_3;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_3;
  wire p_isFull_Pushing_data_to_full_FIFO_prb_4;
  wire p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_4;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_prb_4;
  wire p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_4;
  wire and_244_nl;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_prb_4;
  wire p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_4;
  wire mux_4_nl;
  wire mux_nl;
  wire or_618_nl;
  wire nand_nl;
  wire nor_88_nl;
  wire regIn_chan_TransferNBWrite_if_if_or_nl;
  wire[2:0] regIn_chan_TransferNBWrite_if_if_mux1h_3_nl;
  wire and_nl;
  wire or_590_nl;
  wire[15:0] while_if_for_1_for_acc_nl;
  wire[16:0] nl_while_if_for_1_for_acc_nl;
  wire[15:0] while_if_for_1_for_mux_44_nl;
  wire[15:0] while_if_for_4_and_3_nl;
  wire while_if_for_4_not_2_nl;
  wire or_422_nl;
  wire and_613_nl;
  wire mux_7_nl;
  wire or_635_nl;
  wire or_634_nl;
  wire and_620_nl;
  wire mux_9_nl;
  wire or_639_nl;
  wire nor_90_nl;
  wire and_627_nl;
  wire mux_11_nl;
  wire nand_18_nl;
  wire nor_91_nl;
  wire and_634_nl;
  wire mux_13_nl;
  wire or_648_nl;
  wire or_646_nl;
  wire and_641_nl;
  wire mux_15_nl;
  wire or_653_nl;
  wire or_651_nl;
  wire and_648_nl;
  wire mux_17_nl;
  wire or_656_nl;
  wire nor_94_nl;
  wire and_655_nl;
  wire mux_19_nl;
  wire or_659_nl;
  wire nor_96_nl;
  wire and_662_nl;
  wire mux_21_nl;
  wire or_662_nl;
  wire nor_97_nl;
  wire and_669_nl;
  wire mux_23_nl;
  wire or_666_nl;
  wire or_665_nl;
  wire and_676_nl;
  wire mux_25_nl;
  wire or_670_nl;
  wire or_669_nl;
  wire and_683_nl;
  wire mux_27_nl;
  wire or_673_nl;
  wire nor_98_nl;
  wire and_690_nl;
  wire mux_29_nl;
  wire nand_22_nl;
  wire nor_99_nl;
  wire and_697_nl;
  wire mux_31_nl;
  wire or_681_nl;
  wire or_679_nl;
  wire and_704_nl;
  wire mux_33_nl;
  wire or_686_nl;
  wire or_684_nl;
  wire while_if_for_1_while_if_for_1_nand_2_nl;
  wire and_711_nl;
  wire while_if_for_1_while_if_for_1_nand_1_nl;
  wire and_718_nl;
  wire and_725_nl;
  wire in_or_14_nl;
  wire[15:0] while_if_for_4_and_4_nl;
  wire while_if_for_4_not_3_nl;
  wire or_534_nl;
  wire[15:0] while_if_for_4_and_5_nl;
  wire while_if_for_4_not_4_nl;
  wire or_543_nl;
  wire[1:0] while_if_for_for_b_while_if_for_for_b_mux_nl;
  wire nor_62_nl;
  wire regwr_data_not_nl;
  wire[15:0] mux1h_nl;
  wire and_806_nl;
  wire or_558_nl;
  wire nor_61_nl;
  wire mux_40_nl;
  wire mux_39_nl;
  wire mux_38_nl;
  wire mux_37_nl;
  wire or_718_nl;
  wire mux_35_nl;
  wire axi_read_ar_read_reset_check_ResetChecker_mux_nl;
  wire while_if_for_2_for_while_if_for_2_for_or_nl;
  wire[4:0] while_if_for_1_for_1_acc_1_nl;
  wire[5:0] nl_while_if_for_1_for_1_acc_1_nl;
  wire[3:0] while_if_for_2_for_nor_nl;
  wire in_and_nl;
  wire in_and_1_nl;
  wire in_and_2_nl;
  wire in_and_3_nl;
  wire in_and_4_nl;
  wire in_and_5_nl;
  wire in_and_6_nl;
  wire in_and_7_nl;
  wire in_and_8_nl;
  wire in_and_9_nl;
  wire in_and_10_nl;
  wire in_and_11_nl;
  wire in_and_12_nl;
  wire in_and_13_nl;
  wire in_and_14_nl;
  wire in_and_15_nl;
  wire[3:0] while_if_for_1_for_m_while_if_for_1_for_m_and_nl;
  wire or_573_nl;
  wire and_846_nl;
  wire and_853_nl;
  wire and_860_nl;
  wire operator_64_false_and_2_nl;
  wire operator_64_false_and_3_nl;
  wire operator_64_false_and_4_nl;
  wire operator_64_false_and_5_nl;
  wire operator_64_false_and_10_nl;
  wire operator_64_false_and_11_nl;
  wire operator_64_false_and_12_nl;
  wire operator_64_false_and_13_nl;
  wire operator_64_false_and_18_nl;
  wire operator_64_false_and_19_nl;
  wire operator_64_false_and_20_nl;
  wire operator_64_false_and_21_nl;
  wire operator_64_false_and_26_nl;
  wire operator_64_false_and_27_nl;
  wire operator_64_false_and_28_nl;
  wire operator_64_false_and_29_nl;
  wire[15:0] while_if_for_1_for_mux_39_nl;
  wire[15:0] while_if_for_1_for_mux_41_nl;
  wire[1:0] while_if_for_1_for_while_if_for_1_for_and_1_nl;
  wire while_if_for_1_for_nor_1_nl;
  wire[1:0] while_if_for_1_for_mux1h_1_nl;
  wire while_if_for_1_for_or_1_nl;
  wire[1:0] while_if_for_4_for_mux_39_nl;
  wire or_719_nl;

  // Interconnect Declarations for Component Instantiations 
  wire while_if_for_1_or_nl;
  wire [15:0] nl_while_if_for_1_lshift_rg_a;
  assign while_if_for_1_or_nl = (fsm_output[18]) | (fsm_output[23]);
  assign nl_while_if_for_1_lshift_rg_a = MUX1HOT_v_16_3_2(while_if_for_1_for_mux_38,
      while_if_for_2_for_while_if_for_2_for_mux_2, z_out_4, {(fsm_output[8]) , (fsm_output[13])
      , while_if_for_1_or_nl});
  wire [5:0] nl_while_if_for_1_lshift_rg_s;
  assign nl_while_if_for_1_lshift_rg_s = {while_if_for_1_j_2_0_sva_1_0 , 4'b0000};
  wire  nl_Accelerator_run_run_run_fsm_inst_while_C_1_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_C_1_tr0 = ~ while_lor_lpi_1_dfm_st;
  wire  nl_Accelerator_run_run_run_fsm_inst_while_if_for_for_C_0_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_if_for_for_C_0_tr0 = z_out[2];
  wire  nl_Accelerator_run_run_run_fsm_inst_while_if_for_C_0_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_if_for_C_0_tr0 = z_out[2];
  wire  nl_Accelerator_run_run_run_fsm_inst_while_if_for_1_C_1_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_if_for_1_C_1_tr0 = z_out[2];
  wire  nl_Accelerator_run_run_run_fsm_inst_while_C_2_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_C_2_tr0 = ~ while_lor_lpi_1_dfm_st;
  wire  nl_Accelerator_run_run_run_fsm_inst_while_if_for_2_C_1_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_if_for_2_C_1_tr0 = z_out[2];
  wire  nl_Accelerator_run_run_run_fsm_inst_while_C_3_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_C_3_tr0 = ~ while_lor_lpi_1_dfm_st;
  wire  nl_Accelerator_run_run_run_fsm_inst_while_if_for_3_C_1_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_if_for_3_C_1_tr0 = z_out[2];
  wire  nl_Accelerator_run_run_run_fsm_inst_while_C_4_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_C_4_tr0 = ~ while_lor_lpi_1_dfm_st;
  wire  nl_Accelerator_run_run_run_fsm_inst_while_if_for_4_C_1_tr0;
  assign nl_Accelerator_run_run_run_fsm_inst_while_if_for_4_C_1_tr0 = while_if_for_4_acc_1_cse_1_sva[2];
  mgc_shift_l_v5 #(.width_a(32'sd16),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd64)) while_if_for_1_lshift_rg (
      .a(nl_while_if_for_1_lshift_rg_a[15:0]),
      .s(nl_while_if_for_1_lshift_rg_s[5:0]),
      .z(z_out_3)
    );
  Accelerator_run_run_run_fsm Accelerator_run_run_run_fsm_inst (
      .clk(clk),
      .reset_bar(reset_bar),
      .fsm_output(fsm_output),
      .while_C_1_tr0(nl_Accelerator_run_run_run_fsm_inst_while_C_1_tr0),
      .while_if_for_for_C_0_tr0(nl_Accelerator_run_run_run_fsm_inst_while_if_for_for_C_0_tr0),
      .while_if_for_C_0_tr0(nl_Accelerator_run_run_run_fsm_inst_while_if_for_C_0_tr0),
      .while_if_for_1_for_C_1_tr0(and_dcpl_37),
      .while_if_for_1_C_1_tr0(nl_Accelerator_run_run_run_fsm_inst_while_if_for_1_C_1_tr0),
      .while_C_2_tr0(nl_Accelerator_run_run_run_fsm_inst_while_C_2_tr0),
      .while_if_for_2_for_C_1_tr0(and_dcpl_37),
      .while_if_for_2_C_1_tr0(nl_Accelerator_run_run_run_fsm_inst_while_if_for_2_C_1_tr0),
      .while_C_3_tr0(nl_Accelerator_run_run_run_fsm_inst_while_C_3_tr0),
      .while_if_for_3_for_C_1_tr0(and_dcpl_37),
      .while_if_for_3_C_1_tr0(nl_Accelerator_run_run_run_fsm_inst_while_if_for_3_C_1_tr0),
      .while_C_4_tr0(nl_Accelerator_run_run_run_fsm_inst_while_C_4_tr0),
      .while_if_for_4_for_C_1_tr0(and_dcpl_37),
      .while_if_for_4_C_1_tr0(nl_Accelerator_run_run_run_fsm_inst_while_if_for_4_C_1_tr0)
    );
  assign or_165_cse = mux_1_cse & (regOut_chan_1[2]) & (fsm_output[1]);
  assign p_isFull_Pushing_data_to_full_FIFO_prb = MUX1HOT_s_1_1_2(~ regIn_chan_fifo_write_valid_1_sva,
      or_165_cse);
  // assert(!isFull() && "Pushing data to full FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 247
  property Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isFull_Pushing_data_to_full_FIFO_ctrl_prb  |-> p_isFull_Pushing_data_to_full_FIFO_prb );
  endproperty
  Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO: assert property (Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_p);

  assign regIn_chan_fifo_write_push_mux_1_cse = MUX1HOT_s_1_1_2(1'b1, or_165_cse);
  assign p_isFull_Pushing_data_to_full_FIFO_ctrl_prb = regIn_chan_fifo_write_push_mux_1_cse;
  assign p_isEmpty_Peeking_data_from_empty_FIFO_prb = regIn_chan_fifo_write_push_mux_1_cse;
  // assert(!isEmpty() && "Peeking data from empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 266
  property Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb  |-> p_isEmpty_Peeking_data_from_empty_FIFO_prb );
  endproperty
  Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO: assert property (Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_p);

  assign p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb = regIn_chan_fifo_write_push_mux_1_cse;
  assign and_104_nl = and_dcpl_1 & (fsm_output[2]);
  assign regIn_chan_fifo_write_incrHead_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_104_nl);
  assign p_isEmpty_Incrementing_head_of_empty_FIFO_prb = regIn_chan_fifo_write_incrHead_mux_cse;
  // assert(!isEmpty() && "Incrementing head of empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 260
  property Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb  |-> p_isEmpty_Incrementing_head_of_empty_FIFO_prb );
  endproperty
  Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO: assert property (Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_p);

  assign p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb = regIn_chan_fifo_write_incrHead_mux_cse;
  assign p_isFull_Pushing_data_to_full_FIFO_prb_1 = MUX1HOT_s_1_1_2(regIn_chan_TransferNBWrite_1_if_asn_mdf_sva,
      and_189_cse);
  // assert(!isFull() && "Pushing data to full FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 247
  property Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_1_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_1  |-> p_isFull_Pushing_data_to_full_FIFO_prb_1 );
  endproperty
  Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_1: assert property (Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_1_p);

  assign regIn_chan_fifo_write_push_1_mux_1_cse = MUX1HOT_s_1_1_2(1'b1, and_189_cse);
  assign p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_1 = regIn_chan_fifo_write_push_1_mux_1_cse;
  assign p_isEmpty_Peeking_data_from_empty_FIFO_prb_1 = regIn_chan_fifo_write_push_1_mux_1_cse;
  // assert(!isEmpty() && "Peeking data from empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 266
  property Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_1_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_1  |-> p_isEmpty_Peeking_data_from_empty_FIFO_prb_1 );
  endproperty
  Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_1: assert property (Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_1_p);

  assign p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_1 = regIn_chan_fifo_write_push_1_mux_1_cse;
  assign and_217_nl = and_dcpl_1 & (fsm_output[9]);
  assign regIn_chan_fifo_write_incrHead_1_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_217_nl);
  assign p_isEmpty_Incrementing_head_of_empty_FIFO_prb_1 = regIn_chan_fifo_write_incrHead_1_mux_cse;
  // assert(!isEmpty() && "Incrementing head of empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 260
  property Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_1_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_1  |-> p_isEmpty_Incrementing_head_of_empty_FIFO_prb_1 );
  endproperty
  Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_1: assert property (Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_1_p);

  assign p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_1 = regIn_chan_fifo_write_incrHead_1_mux_cse;
  assign p_isFull_Pushing_data_to_full_FIFO_prb_2 = MUX1HOT_s_1_1_2(regIn_chan_TransferNBWrite_1_if_asn_mdf_sva,
      and_219_cse);
  // assert(!isFull() && "Pushing data to full FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 247
  property Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_2_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_2  |-> p_isFull_Pushing_data_to_full_FIFO_prb_2 );
  endproperty
  Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_2: assert property (Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_2_p);

  assign regIn_chan_fifo_write_push_2_mux_1_cse = MUX1HOT_s_1_1_2(1'b1, and_219_cse);
  assign p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_2 = regIn_chan_fifo_write_push_2_mux_1_cse;
  assign p_isEmpty_Peeking_data_from_empty_FIFO_prb_2 = regIn_chan_fifo_write_push_2_mux_1_cse;
  // assert(!isEmpty() && "Peeking data from empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 266
  property Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_2_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_2  |-> p_isEmpty_Peeking_data_from_empty_FIFO_prb_2 );
  endproperty
  Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_2: assert property (Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_2_p);

  assign p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_2 = regIn_chan_fifo_write_push_2_mux_1_cse;
  assign and_223_nl = and_dcpl_1 & (fsm_output[14]);
  assign regIn_chan_fifo_write_incrHead_2_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_223_nl);
  assign p_isEmpty_Incrementing_head_of_empty_FIFO_prb_2 = regIn_chan_fifo_write_incrHead_2_mux_cse;
  // assert(!isEmpty() && "Incrementing head of empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 260
  property Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_2_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_2  |-> p_isEmpty_Incrementing_head_of_empty_FIFO_prb_2 );
  endproperty
  Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_2: assert property (Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_2_p);

  assign p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_2 = regIn_chan_fifo_write_incrHead_2_mux_cse;
  assign p_isFull_Pushing_data_to_full_FIFO_prb_3 = MUX1HOT_s_1_1_2(regIn_chan_TransferNBWrite_1_if_asn_mdf_sva,
      and_225_cse);
  // assert(!isFull() && "Pushing data to full FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 247
  property Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_3_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_3  |-> p_isFull_Pushing_data_to_full_FIFO_prb_3 );
  endproperty
  Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_3: assert property (Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_3_p);

  assign regIn_chan_fifo_write_push_3_mux_1_cse = MUX1HOT_s_1_1_2(1'b1, and_225_cse);
  assign p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_3 = regIn_chan_fifo_write_push_3_mux_1_cse;
  assign p_isEmpty_Peeking_data_from_empty_FIFO_prb_3 = regIn_chan_fifo_write_push_3_mux_1_cse;
  // assert(!isEmpty() && "Peeking data from empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 266
  property Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_3_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_3  |-> p_isEmpty_Peeking_data_from_empty_FIFO_prb_3 );
  endproperty
  Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_3: assert property (Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_3_p);

  assign p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_3 = regIn_chan_fifo_write_push_3_mux_1_cse;
  assign and_229_nl = and_dcpl_1 & (fsm_output[19]);
  assign regIn_chan_fifo_write_incrHead_3_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_229_nl);
  assign p_isEmpty_Incrementing_head_of_empty_FIFO_prb_3 = regIn_chan_fifo_write_incrHead_3_mux_cse;
  // assert(!isEmpty() && "Incrementing head of empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 260
  property Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_3_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_3  |-> p_isEmpty_Incrementing_head_of_empty_FIFO_prb_3 );
  endproperty
  Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_3: assert property (Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_3_p);

  assign p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_3 = regIn_chan_fifo_write_incrHead_3_mux_cse;
  assign p_isFull_Pushing_data_to_full_FIFO_prb_4 = MUX1HOT_s_1_1_2(regIn_chan_TransferNBWrite_1_if_asn_mdf_sva,
      and_919_cse);
  // assert(!isFull() && "Pushing data to full FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 247
  property Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_4_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_4  |-> p_isFull_Pushing_data_to_full_FIFO_prb_4 );
  endproperty
  Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_4: assert property (Accelerator_run_fifo_h_ln247_assert_not_isFullOP_CP_and_PushingdatatofullFIFO_4_p);

  assign regIn_chan_fifo_write_push_4_mux_1_cse = MUX1HOT_s_1_1_2(1'b1, and_919_cse);
  assign p_isFull_Pushing_data_to_full_FIFO_ctrl_prb_4 = regIn_chan_fifo_write_push_4_mux_1_cse;
  assign p_isEmpty_Peeking_data_from_empty_FIFO_prb_4 = regIn_chan_fifo_write_push_4_mux_1_cse;
  // assert(!isEmpty() && "Peeking data from empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 266
  property Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_4_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_4  |-> p_isEmpty_Peeking_data_from_empty_FIFO_prb_4 );
  endproperty
  Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_4: assert property (Accelerator_run_fifo_h_ln266_assert_not_isEmptyOP_CP_and_PeekingdatafromemptyFIFO_4_p);

  assign p_isEmpty_Peeking_data_from_empty_FIFO_ctrl_prb_4 = regIn_chan_fifo_write_push_4_mux_1_cse;
  assign and_244_nl = and_dcpl_1 & (fsm_output[24]);
  assign regIn_chan_fifo_write_incrHead_4_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_244_nl);
  assign p_isEmpty_Incrementing_head_of_empty_FIFO_prb_4 = regIn_chan_fifo_write_incrHead_4_mux_cse;
  // assert(!isEmpty() && "Incrementing head of empty FIFO") - /mnt/coe/workspace/ece/ece720-common/tools/2020.05/matchlib/cmod/include/fifo.h: line 260
  property Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_4_p;
    @(posedge clk) disable iff ( !reset_bar )
    ( p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_4  |-> p_isEmpty_Incrementing_head_of_empty_FIFO_prb_4 );
  endproperty
  Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_4: assert property (Accelerator_run_fifo_h_ln260_assert_not_isEmptyOP_CP_and_IncrementingheadofemptyFIFO_4_p);

  assign p_isEmpty_Incrementing_head_of_empty_FIFO_ctrl_prb_4 = regIn_chan_fifo_write_incrHead_4_mux_cse;
  assign and_919_cse = (while_if_for_4_acc_1_cse_1_sva[2]) & (fsm_output[23]);
  assign or_618_nl = (regOut_chan_1[0]) | and_tmp;
  assign nand_nl = ~((regOut_chan_1[0]) & (~ and_tmp));
  assign mux_nl = MUX_s_1_2_2(or_618_nl, nand_nl, regOut_chan_1[1]);
  assign nor_88_nl = ~((regOut_chan_1[63:2]!=62'b00000000000000000000000000000000000000000000000000000000000001)
      | (~ (fsm_output[1])));
  assign mux_4_nl = MUX_s_1_2_2(and_tmp, mux_nl, nor_88_nl);
  assign or_619_cse = mux_4_nl | and_919_cse;
  assign regIn_chan_PushNB_mioi_idat = {reg_regIn_chan_PushNB_mioi_idat_ftd , reg_regIn_chan_PushNB_mioi_idat_1_ftd_3
      , reg_regIn_chan_PushNB_mioi_idat_1_ftd_2_0 , 3'b000};
  assign and_nl = (~((regOut_chan_1[63:3]!=61'b0000000000000000000000000000000000000000000000000000000000000)))
      & (regOut_chan_1[0]);
  assign or_590_nl = operator_64_false_1_nor_tmp | (while_if_nor_1_tmp & (regOut_chan_1[0]));
  assign mux_1_cse = MUX_s_1_2_2(and_nl, or_590_nl, regOut_chan_1[1]);
  assign and_107_cse = and_dcpl_3 & (~ (fsm_output[1]));
  assign out_or_cse = (fsm_output[6]) | (fsm_output[11]);
  assign and_508_cse = while_if_for_4_and_tmp_2_sva & (fsm_output[22]);
  assign or_629_cse = (fsm_output[17]) | (fsm_output[15]);
  assign or_636_cse = (fsm_output[0]) | (fsm_output[24]) | (fsm_output[1]) | (fsm_output[2]);
  assign or_633_cse = (fsm_output[6]) | (fsm_output[11]) | (fsm_output[16]) | (fsm_output[21]);
  assign nand_19_cse = ~((while_if_for_2_for_1_acc_1_tmp[3:2]==2'b11));
  assign while_if_for_1_while_if_for_1_nand_2_nl = ~((while_if_for_1_j_2_0_sva_1_0==2'b01));
  assign while_if_for_1_and_5_cse = MUX_v_16_2_2(16'b0000000000000000, out_1_lpi_2,
      while_if_for_1_while_if_for_1_nand_2_nl);
  assign while_if_for_1_while_if_for_1_nand_1_nl = ~((while_if_for_1_j_2_0_sva_1_0==2'b10));
  assign while_if_for_1_and_4_cse = MUX_v_16_2_2(16'b0000000000000000, out_10_lpi_2,
      while_if_for_1_while_if_for_1_nand_1_nl);
  assign and_753_cse = while_if_for_4_and_tmp_1_sva & (fsm_output[22]);
  assign nand_11_cse = ~((while_if_for_1_j_2_0_sva_1_0==2'b11));
  assign and_774_cse = while_if_for_4_and_tmp_sva & (fsm_output[22]);
  assign while_if_for_1_while_if_for_1_or_1_cse = (while_if_for_1_j_2_0_sva_1_0!=2'b00);
  assign or_716_cse = (fsm_output[15]) | (fsm_output[5]) | (fsm_output[10]);
  assign and_809_cse = (while_if_for_4_acc_1_cse_1_sva[2]) & (fsm_output[22]);
  assign in_equal_cse = ~((while_if_for_1_j_2_0_sva_1_0!=2'b00));
  assign in_equal_1_cse = (while_if_for_1_j_2_0_sva_1_0==2'b01);
  assign in_equal_2_cse = (while_if_for_1_j_2_0_sva_1_0==2'b10);
  assign in_equal_3_cse = (while_if_for_1_j_2_0_sva_1_0==2'b11);
  assign while_if_for_1_for_m_while_if_for_1_for_m_and_nl = MUX_v_4_2_2(4'b0000,
      while_if_for_1_for_m_4_0_sva_1_3_0, or_tmp_333);
  assign or_573_nl = or_dcpl_55 | (fsm_output[15]) | (fsm_output[7]) | or_dcpl_209
      | (fsm_output[20]) | (fsm_output[22]);
  assign while_if_for_1_for_m_mux_1_rgt = MUX_v_5_2_2(z_out, ({1'b0 , while_if_for_1_for_m_while_if_for_1_for_m_and_nl}),
      or_573_nl);
  assign nor_104_cse = ~((fsm_output[17]) | (fsm_output[12]));
  assign operator_64_false_1_nor_tmp = ~((regOut_chan_1[63]) | (regOut_chan_1[62])
      | (regOut_chan_1[61]) | (regOut_chan_1[60]) | (regOut_chan_1[59]) | (regOut_chan_1[58])
      | (regOut_chan_1[57]) | (regOut_chan_1[56]) | (regOut_chan_1[55]) | (regOut_chan_1[54])
      | (regOut_chan_1[53]) | (regOut_chan_1[52]) | (regOut_chan_1[51]) | (regOut_chan_1[50])
      | (regOut_chan_1[49]) | (regOut_chan_1[48]) | (regOut_chan_1[47]) | (regOut_chan_1[46])
      | (regOut_chan_1[45]) | (regOut_chan_1[44]) | (regOut_chan_1[43]) | (regOut_chan_1[42])
      | (regOut_chan_1[41]) | (regOut_chan_1[40]) | (regOut_chan_1[39]) | (regOut_chan_1[38])
      | (regOut_chan_1[37]) | (regOut_chan_1[36]) | (regOut_chan_1[35]) | (regOut_chan_1[34])
      | (regOut_chan_1[33]) | (regOut_chan_1[32]) | (regOut_chan_1[31]) | (regOut_chan_1[30])
      | (regOut_chan_1[29]) | (regOut_chan_1[28]) | (regOut_chan_1[27]) | (regOut_chan_1[26])
      | (regOut_chan_1[25]) | (regOut_chan_1[24]) | (regOut_chan_1[23]) | (regOut_chan_1[22])
      | (regOut_chan_1[21]) | (regOut_chan_1[20]) | (regOut_chan_1[19]) | (regOut_chan_1[18])
      | (regOut_chan_1[17]) | (regOut_chan_1[16]) | (regOut_chan_1[15]) | (regOut_chan_1[14])
      | (regOut_chan_1[13]) | (regOut_chan_1[12]) | (regOut_chan_1[11]) | (regOut_chan_1[10])
      | (regOut_chan_1[9]) | (regOut_chan_1[8]) | (regOut_chan_1[7]) | (regOut_chan_1[6])
      | (regOut_chan_1[5]) | (regOut_chan_1[4]) | (regOut_chan_1[3]) | (regOut_chan_1[0]));
  assign while_if_nor_1_tmp = ~((regOut_chan_1[63]) | (regOut_chan_1[62]) | (regOut_chan_1[61])
      | (regOut_chan_1[60]) | (regOut_chan_1[59]) | (regOut_chan_1[58]) | (regOut_chan_1[57])
      | (regOut_chan_1[56]) | (regOut_chan_1[55]) | (regOut_chan_1[54]) | (regOut_chan_1[53])
      | (regOut_chan_1[52]) | (regOut_chan_1[51]) | (regOut_chan_1[50]) | (regOut_chan_1[49])
      | (regOut_chan_1[48]) | (regOut_chan_1[47]) | (regOut_chan_1[46]) | (regOut_chan_1[45])
      | (regOut_chan_1[44]) | (regOut_chan_1[43]) | (regOut_chan_1[42]) | (regOut_chan_1[41])
      | (regOut_chan_1[40]) | (regOut_chan_1[39]) | (regOut_chan_1[38]) | (regOut_chan_1[37])
      | (regOut_chan_1[36]) | (regOut_chan_1[35]) | (regOut_chan_1[34]) | (regOut_chan_1[33])
      | (regOut_chan_1[32]) | (regOut_chan_1[31]) | (regOut_chan_1[30]) | (regOut_chan_1[29])
      | (regOut_chan_1[28]) | (regOut_chan_1[27]) | (regOut_chan_1[26]) | (regOut_chan_1[25])
      | (regOut_chan_1[24]) | (regOut_chan_1[23]) | (regOut_chan_1[22]) | (regOut_chan_1[21])
      | (regOut_chan_1[20]) | (regOut_chan_1[19]) | (regOut_chan_1[18]) | (regOut_chan_1[17])
      | (regOut_chan_1[16]) | (regOut_chan_1[15]) | (regOut_chan_1[14]) | (regOut_chan_1[13])
      | (regOut_chan_1[12]) | (regOut_chan_1[11]) | (regOut_chan_1[10]) | (regOut_chan_1[9])
      | (regOut_chan_1[8]) | (regOut_chan_1[7]) | (regOut_chan_1[6]) | (regOut_chan_1[5])
      | (regOut_chan_1[4]) | (regOut_chan_1[3]) | (regOut_chan_1[1]));
  assign out_3_sva_1_mx0w0 = MUX_v_16_2_2(16'b0000000000000000, out_11_lpi_2, nand_11_cse);
  assign operator_64_false_and_2_nl = in_equal_cse & operator_64_false_nor_m1c_1;
  assign operator_64_false_and_3_nl = in_equal_1_cse & operator_64_false_nor_m1c_1;
  assign operator_64_false_and_4_nl = in_equal_2_cse & operator_64_false_nor_m1c_1;
  assign operator_64_false_and_5_nl = in_equal_3_cse & operator_64_false_nor_m1c_1;
  assign operator_64_false_and_10_nl = in_equal_cse & operator_64_false_and_m1c_3;
  assign operator_64_false_and_11_nl = in_equal_1_cse & operator_64_false_and_m1c_3;
  assign operator_64_false_and_12_nl = in_equal_2_cse & operator_64_false_and_m1c_3;
  assign operator_64_false_and_13_nl = in_equal_3_cse & operator_64_false_and_m1c_3;
  assign operator_64_false_and_18_nl = in_equal_cse & operator_64_false_and_m1c_4;
  assign operator_64_false_and_19_nl = in_equal_1_cse & operator_64_false_and_m1c_4;
  assign operator_64_false_and_20_nl = in_equal_2_cse & operator_64_false_and_m1c_4;
  assign operator_64_false_and_21_nl = in_equal_3_cse & operator_64_false_and_m1c_4;
  assign operator_64_false_and_26_nl = in_equal_cse & operator_64_false_and_m1c_5;
  assign operator_64_false_and_27_nl = in_equal_1_cse & operator_64_false_and_m1c_5;
  assign operator_64_false_and_28_nl = in_equal_2_cse & operator_64_false_and_m1c_5;
  assign operator_64_false_and_29_nl = in_equal_3_cse & operator_64_false_and_m1c_5;
  assign operator_64_false_rshift_ctmp_sva_2 = MUX1HOT_v_16_16_2((regOut_chan_2[15:0]),
      (regOut_chan_3[15:0]), (regOut_chan_4[15:0]), (regOut_chan_5[15:0]), (regOut_chan_2[31:16]),
      (regOut_chan_3[31:16]), (regOut_chan_4[31:16]), (regOut_chan_5[31:16]), (regOut_chan_2[47:32]),
      (regOut_chan_3[47:32]), (regOut_chan_4[47:32]), (regOut_chan_5[47:32]), (regOut_chan_2[63:48]),
      (regOut_chan_3[63:48]), (regOut_chan_4[63:48]), (regOut_chan_5[63:48]), {operator_64_false_and_2_nl
      , operator_64_false_and_3_nl , operator_64_false_and_4_nl , operator_64_false_and_5_nl
      , operator_64_false_and_10_nl , operator_64_false_and_11_nl , operator_64_false_and_12_nl
      , operator_64_false_and_13_nl , operator_64_false_and_18_nl , operator_64_false_and_19_nl
      , operator_64_false_and_20_nl , operator_64_false_and_21_nl , operator_64_false_and_26_nl
      , operator_64_false_and_27_nl , operator_64_false_and_28_nl , operator_64_false_and_29_nl});
  assign operator_64_false_nor_m1c_1 = ~((while_if_for_for_b_2_0_sva_1_0!=2'b00));
  assign operator_64_false_and_m1c_3 = (while_if_for_for_b_2_0_sva_1_0==2'b01);
  assign operator_64_false_and_m1c_4 = (while_if_for_for_b_2_0_sva_1_0==2'b10);
  assign operator_64_false_and_m1c_5 = (while_if_for_for_b_2_0_sva_1_0==2'b11);
  assign regwr_data_1_sva_2 = regwr_data_1_sva | z_out_3;
  assign while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1 =
      MUX_v_16_16_2x0(in_1_lpi_3, in_2_lpi_3, in_3_lpi_3, in_4_lpi_3, in_5_lpi_3,
      in_6_lpi_3, in_7_lpi_3, in_8_lpi_3, in_9_lpi_3, in_10_lpi_3, in_11_lpi_3, in_12_lpi_3,
      in_13_lpi_3, in_14_lpi_3, in_15_1_sva, while_if_for_2_for_1_acc_1_tmp);
  assign nl_while_if_for_2_for_1_acc_1_tmp = while_if_for_1_for_1_n_3_0_sva + 4'b0001;
  assign while_if_for_2_for_1_acc_1_tmp = nl_while_if_for_2_for_1_acc_1_tmp[3:0];
  assign while_if_for_4_and_tmp_sva_mx0w0 = (z_out[1:0]==2'b11);
  assign while_if_for_4_and_tmp_1_sva_mx0w0 = (z_out[1:0]==2'b10);
  assign while_if_for_4_and_tmp_2_sva_mx0w0 = (z_out[1:0]==2'b01);
  assign while_if_for_1_for_mux_38 = MUX_v_16_4_2(out_0_lpi_2, out_1_sva_1, out_2_sva_1,
      out_3_sva_1, while_if_for_1_j_2_0_sva_1_0);
  assign while_if_for_2_for_while_if_for_2_for_mux_2 = MUX_v_16_4_2(out_0_lpi_2,
      out_5_sva_1, out_6_sva_1, out_7_sva_1, while_if_for_1_j_2_0_sva_1_0);
  assign while_if_for_1_for_mux_39_nl = MUX_v_16_16_2(we_0_lpi_3, we_1_lpi_3, we_2_lpi_3,
      we_3_lpi_3, we_4_lpi_3, we_5_lpi_3, we_6_lpi_3, we_7_lpi_3, we_8_lpi_3, we_9_lpi_3,
      we_10_lpi_3, we_11_lpi_3, we_12_lpi_3, we_13_lpi_3, we_14_lpi_3, we_15_lpi_3,
      while_if_for_1_for_m_4_0_sva_1_3_0);
  assign while_if_for_1_for_mux_41_nl = MUX_v_16_16_2(in_0_lpi_3, in_1_lpi_3, in_2_lpi_3,
      in_3_lpi_3, in_4_lpi_3, in_5_lpi_3, in_6_lpi_3, in_7_lpi_3, in_8_lpi_3, in_9_lpi_3,
      in_10_lpi_3, in_11_lpi_3, in_12_lpi_3, in_13_lpi_3, in_14_lpi_3, in_15_1_sva,
      while_if_for_1_for_m_4_0_sva_1_3_0);
  assign nl_while_if_for_1_for_mul_2 = $signed(while_if_for_1_for_mux_39_nl) * $signed(while_if_for_1_for_mux_41_nl);
  assign while_if_for_1_for_mul_2 = nl_while_if_for_1_for_mul_2[15:0];
  assign and_dcpl_1 = while_lor_lpi_1_dfm_st & regIn_chan_PushNB_mioi_irdy;
  assign and_dcpl_3 = ~((fsm_output[24]) | (fsm_output[0]));
  assign or_dcpl_55 = (fsm_output[5]) | (fsm_output[10]);
  assign and_189_cse = (z_out[2]) & (fsm_output[8]);
  assign and_219_cse = (z_out[2]) & (fsm_output[13]);
  assign and_225_cse = (z_out[2]) & (fsm_output[18]);
  assign and_dcpl_37 = exit_while_if_for_1_for_1_sva & while_if_for_1_for_m_4_0_sva_1_4;
  assign or_dcpl_135 = (while_if_for_1_j_2_0_sva_1_0!=2'b01);
  assign or_dcpl_136 = ~((while_if_for_for_b_2_0_sva_1_0==2'b11));
  assign or_dcpl_139 = (while_if_for_for_b_2_0_sva_1_0!=2'b00);
  assign or_dcpl_142 = (while_if_for_for_b_2_0_sva_1_0!=2'b10);
  assign or_dcpl_144 = (while_if_for_for_b_2_0_sva_1_0!=2'b01);
  assign or_dcpl_150 = (while_if_for_1_j_2_0_sva_1_0!=2'b10);
  assign and_dcpl_55 = ~((fsm_output[24]) | (fsm_output[1]));
  assign and_dcpl_58 = ~((fsm_output[6]) | (fsm_output[11]));
  assign or_dcpl_165 = out_or_cse | (fsm_output[16]) | (fsm_output[21]);
  assign and_dcpl_61 = (while_if_for_1_for_1_n_3_0_sva[1:0]==2'b01);
  assign and_dcpl_62 = ~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva[3]));
  assign and_dcpl_63 = and_dcpl_62 & (~ (while_if_for_1_for_1_n_3_0_sva[2]));
  assign and_dcpl_65 = (while_if_for_1_for_1_n_3_0_sva[1:0]==2'b10);
  assign and_dcpl_66 = (~ exit_while_if_for_1_for_1_sva) & (while_if_for_1_for_1_n_3_0_sva[3]);
  assign and_dcpl_67 = and_dcpl_66 & (~ (while_if_for_1_for_1_n_3_0_sva[2]));
  assign and_dcpl_69 = (while_if_for_1_for_1_n_3_0_sva[1:0]==2'b11);
  assign and_dcpl_71 = ~((while_if_for_1_for_1_n_3_0_sva[1:0]!=2'b00));
  assign and_dcpl_72 = and_dcpl_66 & (while_if_for_1_for_1_n_3_0_sva[2]);
  assign and_dcpl_78 = and_dcpl_62 & (while_if_for_1_for_1_n_3_0_sva[2]);
  assign or_dcpl_204 = (fsm_output[7]) | (fsm_output[12]);
  assign or_dcpl_208 = (fsm_output[22:21]!=2'b00);
  assign or_dcpl_209 = (fsm_output[12]) | (fsm_output[17]);
  assign or_tmp_141 = while_lor_lpi_1_dfm_st & (fsm_output[24]);
  assign or_tmp_197 = and_107_cse & (fsm_output[3:2]==2'b00);
  assign and_707_cse = (~((fsm_output[5]) | (fsm_output[0]))) & and_dcpl_55 & (~((fsm_output[2])
      | (fsm_output[7]))) & (~((fsm_output[4:3]!=2'b00)));
  assign or_tmp_331 = and_dcpl_58 & (~((fsm_output[16]) | (fsm_output[7]))) & nor_104_cse
      & (fsm_output[22:21]==2'b00);
  assign or_tmp_333 = or_dcpl_204 | (fsm_output[17]) | (fsm_output[22]);
  assign and_842_cse = (fsm_output[15]) | (fsm_output[11]) | (fsm_output[16]) | (fsm_output[17])
      | (fsm_output[13]) | (fsm_output[14]) | (fsm_output[18]) | (fsm_output[19])
      | (fsm_output[23]) | (fsm_output[20]) | (fsm_output[21]) | (fsm_output[22]);
  assign regwr_data_1_sva_mx0c0 = (fsm_output[9]) | (fsm_output[14]) | (fsm_output[19])
      | (fsm_output[4]);
  assign or_601_ssc = (fsm_output[18]) | (fsm_output[13]) | (fsm_output[8]) | (fsm_output[4]);
  assign and_tmp = (z_out[2]) & ((fsm_output[8]) | (fsm_output[13]) | (fsm_output[18]));
  assign or_tmp_432 = (~ (fsm_output[20])) | (z_out[2]);
  assign or_tmp_433 = (while_if_for_1_j_2_0_sva_1_0!=2'b00) | (~ or_tmp_432);
  assign mux_tmp_36 = MUX_s_1_2_2(and_809_cse, (z_out[2]), fsm_output[20]);
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_regIn_chan_PushNB_mioi_idat_ftd <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      reg_regIn_chan_PushNB_mioi_idat_1_ftd_3 <= 1'b0;
      reg_regIn_chan_PushNB_mioi_idat_1_ftd_2_0 <= 3'b000;
    end
    else if ( or_619_cse ) begin
      reg_regIn_chan_PushNB_mioi_idat_ftd <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          regwr_data_1_sva_2, regIn_chan_TransferNBWrite_if_if_or_nl);
      reg_regIn_chan_PushNB_mioi_idat_1_ftd_3 <= ~ or_165_cse;
      reg_regIn_chan_PushNB_mioi_idat_1_ftd_2_0 <= ~(MUX_v_3_2_2(regIn_chan_TransferNBWrite_if_if_mux1h_3_nl,
          3'b111, or_165_cse));
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regIn_chan_PushNB_mioi_ivld <= 1'b0;
      while_if_for_for_b_2_0_sva_1_0 <= 2'b00;
      exit_while_if_for_1_for_1_sva <= 1'b0;
      while_if_for_1_for_m_4_0_sva_1_4 <= 1'b0;
      while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva <= 16'b0000000000000000;
    end
    else begin
      regIn_chan_PushNB_mioi_ivld <= ~(((~((fsm_output[1]) | (fsm_output[8]) | (fsm_output[13])))
          & (~((fsm_output[18]) | (fsm_output[23])))) | ((~ (while_if_for_4_acc_1_cse_1_sva[2]))
          & (fsm_output[23])) | (~((z_out[2]) | (fsm_output[1]) | (fsm_output[23])))
          | ((~(mux_1_cse & (regOut_chan_1[2]))) & (fsm_output[1])));
      while_if_for_for_b_2_0_sva_1_0 <= MUX_v_2_2_2(2'b00, (z_out[1:0]), (fsm_output[3]));
      exit_while_if_for_1_for_1_sva <= axi_read_ar_read_reset_check_ResetChecker_mux_nl
          & (~ or_tmp_331);
      while_if_for_1_for_m_4_0_sva_1_4 <= while_if_for_1_for_m_mux_1_rgt[4];
      while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva <= nl_while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva[15:0];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regIn_chan_fifo_write_valid_1_sva <= 1'b0;
      out_12_sva <= 16'b0000000000000000;
      out_9_sva <= 16'b0000000000000000;
      out_10_sva <= 16'b0000000000000000;
      out_11_sva <= 16'b0000000000000000;
      out_7_sva <= 16'b0000000000000000;
      out_6_sva <= 16'b0000000000000000;
      out_5_sva <= 16'b0000000000000000;
      we_7_sva <= 16'b0000000000000000;
      we_8_sva <= 16'b0000000000000000;
      we_6_sva <= 16'b0000000000000000;
      we_9_sva <= 16'b0000000000000000;
      we_5_sva <= 16'b0000000000000000;
      we_10_sva <= 16'b0000000000000000;
      we_4_sva <= 16'b0000000000000000;
      we_11_sva <= 16'b0000000000000000;
      we_3_sva <= 16'b0000000000000000;
      we_12_sva <= 16'b0000000000000000;
      we_2_sva <= 16'b0000000000000000;
      we_13_sva <= 16'b0000000000000000;
      we_1_sva <= 16'b0000000000000000;
      we_14_sva <= 16'b0000000000000000;
      we_15_sva <= 16'b0000000000000000;
      out_3_sva <= 16'b0000000000000000;
      out_2_sva <= 16'b0000000000000000;
      out_1_sva <= 16'b0000000000000000;
      in_7_sva <= 16'b0000000000000000;
      in_8_sva <= 16'b0000000000000000;
      in_6_sva <= 16'b0000000000000000;
      in_9_sva <= 16'b0000000000000000;
      in_5_sva <= 16'b0000000000000000;
      in_10_sva <= 16'b0000000000000000;
      in_4_sva <= 16'b0000000000000000;
      in_11_sva <= 16'b0000000000000000;
      in_3_sva <= 16'b0000000000000000;
      in_12_sva <= 16'b0000000000000000;
      in_2_sva <= 16'b0000000000000000;
      in_13_sva <= 16'b0000000000000000;
      in_1_sva <= 16'b0000000000000000;
      in_14_sva <= 16'b0000000000000000;
      in_0_sva <= 16'b0000000000000000;
    end
    else if ( or_tmp_141 ) begin
      regIn_chan_fifo_write_valid_1_sva <= ~ regIn_chan_PushNB_mioi_irdy;
      out_12_sva <= out_0_lpi_2;
      out_9_sva <= out_1_lpi_2;
      out_10_sva <= out_10_lpi_2;
      out_11_sva <= out_11_lpi_2;
      out_7_sva <= out_7_sva_1;
      out_6_sva <= out_6_sva_1;
      out_5_sva <= out_5_sva_1;
      we_7_sva <= we_7_lpi_3;
      we_8_sva <= we_8_lpi_3;
      we_6_sva <= we_6_lpi_3;
      we_9_sva <= we_9_lpi_3;
      we_5_sva <= we_5_lpi_3;
      we_10_sva <= we_10_lpi_3;
      we_4_sva <= we_4_lpi_3;
      we_11_sva <= we_11_lpi_3;
      we_3_sva <= we_3_lpi_3;
      we_12_sva <= we_12_lpi_3;
      we_2_sva <= we_2_lpi_3;
      we_13_sva <= we_13_lpi_3;
      we_1_sva <= we_1_lpi_3;
      we_14_sva <= we_14_lpi_3;
      we_15_sva <= we_15_lpi_3;
      out_3_sva <= out_3_sva_1;
      out_2_sva <= out_2_sva_1;
      out_1_sva <= out_1_sva_1;
      in_7_sva <= in_7_lpi_3;
      in_8_sva <= in_8_lpi_3;
      in_6_sva <= in_6_lpi_3;
      in_9_sva <= in_9_lpi_3;
      in_5_sva <= in_5_lpi_3;
      in_10_sva <= in_10_lpi_3;
      in_4_sva <= in_4_lpi_3;
      in_11_sva <= in_11_lpi_3;
      in_3_sva <= in_3_lpi_3;
      in_12_sva <= in_12_lpi_3;
      in_2_sva <= in_2_lpi_3;
      in_13_sva <= in_13_lpi_3;
      in_1_sva <= in_1_lpi_3;
      in_14_sva <= in_14_lpi_3;
      in_0_sva <= in_0_lpi_3;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_lor_lpi_1_dfm_st <= 1'b0;
    end
    else if ( ~ and_107_cse ) begin
      while_lor_lpi_1_dfm_st <= ((regOut_chan_1[2:1]==2'b11) & operator_64_false_1_nor_tmp)
          | ((regOut_chan_1[2]) & (regOut_chan_1[0]) & while_if_nor_1_tmp);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( ((while_if_for_1_j_2_0_sva_1_0==2'b01) & or_629_cse) | and_508_cse
        | ((z_out[1:0]==2'b01) & (fsm_output[20])) | (fsm_output[6]) | (fsm_output[2])
        | (fsm_output[8]) | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13])
        | (fsm_output[14]) ) begin
      out_1_lpi_2 <= MUX1HOT_v_16_9_2(out_1_sva, while_if_for_1_for_acc_nl, out_1_sva_1,
          out_5_sva, out_5_sva_1, out_9_sva, while_if_for_1_and_5_cse, while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva,
          while_if_for_4_and_3_nl, {(fsm_output[2]) , out_or_cse , (fsm_output[8])
          , (fsm_output[9]) , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[15])
          , or_422_nl , (fsm_output[20])});
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_15_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(nand_11_cse | or_dcpl_136 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_15_lpi_3 <= MUX_v_16_2_2(we_15_sva, operator_64_false_rshift_ctmp_sva_2,
          fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_0_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(while_if_for_1_while_if_for_1_or_1_cse | or_dcpl_139 | or_tmp_197)
        ) begin
      we_0_lpi_3 <= operator_64_false_rshift_ctmp_sva_2;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_14_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(nand_11_cse | or_dcpl_142 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_14_lpi_3 <= MUX_v_16_2_2(we_14_sva, operator_64_false_rshift_ctmp_sva_2,
          fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_1_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(while_if_for_1_while_if_for_1_or_1_cse | or_dcpl_144 | or_tmp_197))
        | (fsm_output[2]) ) begin
      we_1_lpi_3 <= MUX_v_16_2_2(we_1_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_13_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(nand_11_cse | or_dcpl_144 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_13_lpi_3 <= MUX_v_16_2_2(we_13_sva, operator_64_false_rshift_ctmp_sva_2,
          fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_2_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(while_if_for_1_while_if_for_1_or_1_cse | or_dcpl_142 | or_tmp_197))
        | (fsm_output[2]) ) begin
      we_2_lpi_3 <= MUX_v_16_2_2(we_2_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_12_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(nand_11_cse | or_dcpl_139 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_12_lpi_3 <= MUX_v_16_2_2(we_12_sva, operator_64_false_rshift_ctmp_sva_2,
          fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_3_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(while_if_for_1_while_if_for_1_or_1_cse | or_dcpl_136 | or_tmp_197))
        | (fsm_output[2]) ) begin
      we_3_lpi_3 <= MUX_v_16_2_2(we_3_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_11_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_150 | or_dcpl_136 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_11_lpi_3 <= MUX_v_16_2_2(we_11_sva, operator_64_false_rshift_ctmp_sva_2,
          fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_4_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_135 | or_dcpl_139 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_4_lpi_3 <= MUX_v_16_2_2(we_4_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_10_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_150 | or_dcpl_142 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_10_lpi_3 <= MUX_v_16_2_2(we_10_sva, operator_64_false_rshift_ctmp_sva_2,
          fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_5_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_135 | or_dcpl_144 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_5_lpi_3 <= MUX_v_16_2_2(we_5_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_9_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_150 | or_dcpl_144 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_9_lpi_3 <= MUX_v_16_2_2(we_9_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_6_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_135 | or_dcpl_142 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_6_lpi_3 <= MUX_v_16_2_2(we_6_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_8_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_150 | or_dcpl_139 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_8_lpi_3 <= MUX_v_16_2_2(we_8_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      we_7_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_135 | or_dcpl_136 | or_tmp_197)) | (fsm_output[2]) ) begin
      we_7_lpi_3 <= MUX_v_16_2_2(we_7_sva, operator_64_false_rshift_ctmp_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regIn_chan_TransferNBWrite_1_if_asn_mdf_sva <= 1'b0;
    end
    else if ( ~(and_dcpl_3 & (~((fsm_output[2:1]!=2'b00))) & (~((fsm_output[9]) |
        (fsm_output[14]))) & (~ (fsm_output[19]))) ) begin
      regIn_chan_TransferNBWrite_1_if_asn_mdf_sva <= regIn_chan_PushNB_mioi_irdy;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_1_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_7_nl, or_633_cse) ) begin
      in_1_lpi_3 <= MUX_v_16_2_2(in_1_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_613_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_10_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_9_nl, or_633_cse) ) begin
      in_10_lpi_3 <= MUX_v_16_2_2(in_10_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_620_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_11_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_11_nl, or_633_cse) ) begin
      in_11_lpi_3 <= MUX_v_16_2_2(in_11_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_627_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_12_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_13_nl, or_633_cse) ) begin
      in_12_lpi_3 <= MUX_v_16_2_2(in_12_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_634_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_13_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_15_nl, or_633_cse) ) begin
      in_13_lpi_3 <= MUX_v_16_2_2(in_13_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_641_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_14_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_17_nl, or_633_cse) ) begin
      in_14_lpi_3 <= MUX_v_16_2_2(in_14_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_648_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_2_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_19_nl, or_633_cse) ) begin
      in_2_lpi_3 <= MUX_v_16_2_2(in_2_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_655_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_3_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_21_nl, or_633_cse) ) begin
      in_3_lpi_3 <= MUX_v_16_2_2(in_3_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_662_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_4_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_23_nl, or_633_cse) ) begin
      in_4_lpi_3 <= MUX_v_16_2_2(in_4_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_669_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_5_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_25_nl, or_633_cse) ) begin
      in_5_lpi_3 <= MUX_v_16_2_2(in_5_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_676_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_6_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_27_nl, or_633_cse) ) begin
      in_6_lpi_3 <= MUX_v_16_2_2(in_6_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_683_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_7_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_29_nl, or_633_cse) ) begin
      in_7_lpi_3 <= MUX_v_16_2_2(in_7_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_690_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_8_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_31_nl, or_633_cse) ) begin
      in_8_lpi_3 <= MUX_v_16_2_2(in_8_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_697_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_9_lpi_3 <= 16'b0000000000000000;
    end
    else if ( MUX_s_1_2_2(or_636_cse, mux_33_nl, or_633_cse) ) begin
      in_9_lpi_3 <= MUX_v_16_2_2(in_9_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          and_704_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_1_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~(and_707_cse | (or_dcpl_135 & (fsm_output[7]))) ) begin
      out_1_sva_1 <= MUX_v_16_2_2(while_if_for_1_and_5_cse, out_1_lpi_2, and_711_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_2_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~(and_707_cse | (or_dcpl_150 & (fsm_output[7]))) ) begin
      out_2_sva_1 <= MUX_v_16_2_2(while_if_for_1_and_4_cse, out_1_lpi_2, and_718_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_3_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~(and_707_cse | (nand_11_cse & (fsm_output[7]))) ) begin
      out_3_sva_1 <= MUX_v_16_2_2(out_3_sva_1_mx0w0, out_1_lpi_2, and_725_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_0_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b0000)
        | (and_dcpl_58 & (~((fsm_output[16]) | (fsm_output[0]))) & and_dcpl_55 &
        (~ (fsm_output[21]))))) | (fsm_output[2]) ) begin
      in_0_lpi_3 <= MUX_v_16_2_2(in_0_sva, while_if_for_1_for_1_while_if_for_1_for_1_slc_in_16_15_0_1_ctmp_sva_1,
          in_or_14_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( ((while_if_for_1_j_2_0_sva_1_0==2'b10) & or_629_cse) | ((z_out[1:0]==2'b10)
        & (fsm_output[20])) | and_753_cse | (fsm_output[2]) | (fsm_output[8]) | (fsm_output[9])
        | (fsm_output[13]) | (fsm_output[14]) ) begin
      out_10_lpi_2 <= MUX1HOT_v_16_8_2(out_2_sva, out_2_sva_1, out_6_sva, out_6_sva_1,
          out_10_sva, while_if_for_1_and_4_cse, while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva,
          while_if_for_4_and_4_nl, {(fsm_output[2]) , (fsm_output[8]) , (fsm_output[9])
          , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[15]) , or_534_nl ,
          (fsm_output[20])});
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( ((while_if_for_1_j_2_0_sva_1_0==2'b11) & or_629_cse) | ((z_out[1:0]==2'b11)
        & (fsm_output[20])) | and_774_cse | (fsm_output[2]) | (fsm_output[8]) | (fsm_output[9])
        | (fsm_output[13]) | (fsm_output[14]) ) begin
      out_11_lpi_2 <= MUX1HOT_v_16_8_2(out_3_sva, out_3_sva_1, out_7_sva, out_7_sva_1,
          out_11_sva, out_3_sva_1_mx0w0, while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva,
          while_if_for_4_and_5_nl, {(fsm_output[2]) , (fsm_output[8]) , (fsm_output[9])
          , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[15]) , or_543_nl ,
          (fsm_output[20])});
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_if_for_1_j_2_0_sva_1_0 <= 2'b00;
    end
    else if ( (fsm_output[23]) | (fsm_output[18]) | (fsm_output[13]) | (fsm_output[8])
        | (fsm_output[4]) | (fsm_output[19]) | (fsm_output[14]) | (fsm_output[2])
        | (fsm_output[9]) ) begin
      while_if_for_1_j_2_0_sva_1_0 <= MUX_v_2_2_2(2'b00, while_if_for_for_b_while_if_for_for_b_mux_nl,
          nor_62_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regwr_data_1_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( regwr_data_1_sva_mx0c0 | (fsm_output[8]) | (fsm_output[13]) | (fsm_output[18])
        | (fsm_output[23]) ) begin
      regwr_data_1_sva <= MUX_v_64_2_2(64'b0000000000000000000000000000000000000000000000000000000000000000,
          regwr_data_1_sva_2, regwr_data_not_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_0_lpi_2 <= 16'b0000000000000000;
    end
    else if ( ~ mux_40_nl ) begin
      out_0_lpi_2 <= MUX_v_16_2_2(16'b0000000000000000, mux1h_nl, nor_61_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_if_for_1_for_1_n_3_0_sva <= 4'b0000;
    end
    else if ( (~((fsm_output[12]) | (fsm_output[7]))) & (~((fsm_output[17]) | (fsm_output[22])))
        ) begin
      while_if_for_1_for_1_n_3_0_sva <= ~(MUX_v_4_2_2(while_if_for_2_for_nor_nl,
          4'b1111, or_tmp_331));
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      in_15_1_sva <= 16'b0000000000000000;
    end
    else if ( ~(out_or_cse | (fsm_output[16]) | (fsm_output[7]) | or_dcpl_209 | or_dcpl_208)
        ) begin
      in_15_1_sva <= MUX1HOT_v_16_16_2((regOut_chan_6[15:0]), (regOut_chan_6[31:16]),
          (regOut_chan_6[47:32]), (regOut_chan_6[63:48]), (regOut_chan_7[15:0]),
          (regOut_chan_7[31:16]), (regOut_chan_7[47:32]), (regOut_chan_7[63:48]),
          (regOut_chan_8[15:0]), (regOut_chan_8[31:16]), (regOut_chan_8[47:32]),
          (regOut_chan_8[63:48]), (regOut_chan_9[15:0]), (regOut_chan_9[31:16]),
          (regOut_chan_9[47:32]), (regOut_chan_9[63:48]), {in_and_nl , in_and_1_nl
          , in_and_2_nl , in_and_3_nl , in_and_4_nl , in_and_5_nl , in_and_6_nl ,
          in_and_7_nl , in_and_8_nl , in_and_9_nl , in_and_10_nl , in_and_11_nl ,
          in_and_12_nl , in_and_13_nl , in_and_14_nl , in_and_15_nl});
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_if_for_1_for_m_4_0_sva_1_3_0 <= 4'b0000;
    end
    else if ( nor_104_cse & (~((fsm_output[7]) | (fsm_output[22]))) ) begin
      while_if_for_1_for_m_4_0_sva_1_3_0 <= while_if_for_1_for_m_mux_1_rgt[3:0];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_5_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~(and_842_cse | (or_dcpl_135 & (fsm_output[12]))) ) begin
      out_5_sva_1 <= MUX_v_16_2_2(while_if_for_1_and_5_cse, out_1_lpi_2, and_846_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_6_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~(and_842_cse | (or_dcpl_150 & (fsm_output[12]))) ) begin
      out_6_sva_1 <= MUX_v_16_2_2(while_if_for_1_and_4_cse, out_1_lpi_2, and_853_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      out_7_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~(and_842_cse | (nand_11_cse & (fsm_output[12]))) ) begin
      out_7_sva_1 <= MUX_v_16_2_2(out_3_sva_1_mx0w0, out_1_lpi_2, and_860_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_if_for_4_acc_1_cse_1_sva <= 3'b000;
    end
    else if ( fsm_output[20] ) begin
      while_if_for_4_acc_1_cse_1_sva <= z_out[2:0];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_if_for_4_and_tmp_sva <= 1'b0;
    end
    else if ( ~ or_dcpl_208 ) begin
      while_if_for_4_and_tmp_sva <= while_if_for_4_and_tmp_sva_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_if_for_4_and_tmp_1_sva <= 1'b0;
    end
    else if ( ~ or_dcpl_208 ) begin
      while_if_for_4_and_tmp_1_sva <= while_if_for_4_and_tmp_1_sva_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_if_for_4_and_tmp_2_sva <= 1'b0;
    end
    else if ( ~ or_dcpl_208 ) begin
      while_if_for_4_and_tmp_2_sva <= while_if_for_4_and_tmp_2_sva_mx0w0;
    end
  end
  assign regIn_chan_TransferNBWrite_if_if_or_nl = and_189_cse | and_219_cse | and_225_cse
      | and_919_cse;
  assign regIn_chan_TransferNBWrite_if_if_mux1h_3_nl = MUX1HOT_v_3_4_2(3'b101, 3'b100,
      3'b011, 3'b010, {and_189_cse , and_219_cse , and_225_cse , and_919_cse});
  assign nl_while_if_for_1_for_1_acc_1_nl = ({1'b1 , while_if_for_2_for_1_acc_1_tmp})
      + 5'b00001;
  assign while_if_for_1_for_1_acc_1_nl = nl_while_if_for_1_for_1_acc_1_nl[4:0];
  assign while_if_for_2_for_while_if_for_2_for_or_nl = (~ (readslicef_5_1_4(while_if_for_1_for_1_acc_1_nl)))
      | exit_while_if_for_1_for_1_sva;
  assign axi_read_ar_read_reset_check_ResetChecker_mux_nl = MUX_s_1_2_2(while_if_for_2_for_while_if_for_2_for_or_nl,
      exit_while_if_for_1_for_1_sva, or_tmp_333);
  assign nl_while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva  = z_out_4 + while_if_for_1_for_mul_2;
  assign while_if_for_1_for_mux_44_nl = MUX_v_16_2_2(while_if_for_1_for_mux_38, while_if_for_2_for_while_if_for_2_for_mux_2,
      fsm_output[11]);
  assign nl_while_if_for_1_for_acc_nl = while_if_for_1_for_mux_44_nl + while_if_for_1_for_mul_2;
  assign while_if_for_1_for_acc_nl = nl_while_if_for_1_for_acc_nl[15:0];
  assign while_if_for_4_not_2_nl = ~ while_if_for_4_and_tmp_2_sva_mx0w0;
  assign while_if_for_4_and_3_nl = MUX_v_16_2_2(16'b0000000000000000, out_1_lpi_2,
      while_if_for_4_not_2_nl);
  assign or_422_nl = (in_equal_1_cse & (fsm_output[17])) | and_508_cse;
  assign and_613_nl = and_dcpl_63 & and_dcpl_61 & or_dcpl_165;
  assign or_635_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b0001);
  assign or_634_nl = exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b0001);
  assign mux_7_nl = MUX_s_1_2_2(or_635_nl, (fsm_output[2]), or_634_nl);
  assign and_620_nl = and_dcpl_67 & and_dcpl_65 & or_dcpl_165;
  assign or_639_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b1010);
  assign nor_90_nl = ~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b1010));
  assign mux_9_nl = MUX_s_1_2_2((fsm_output[2]), or_639_nl, nor_90_nl);
  assign and_627_nl = and_dcpl_67 & and_dcpl_69 & or_dcpl_165;
  assign nand_18_nl = ~((while_if_for_2_for_1_acc_1_tmp==4'b1011));
  assign nor_91_nl = ~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b1011));
  assign mux_11_nl = MUX_s_1_2_2((fsm_output[2]), nand_18_nl, nor_91_nl);
  assign and_634_nl = and_dcpl_72 & and_dcpl_71 & or_dcpl_165;
  assign or_648_nl = (while_if_for_2_for_1_acc_1_tmp[1:0]!=2'b00) | nand_19_cse;
  assign or_646_nl = exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b1100);
  assign mux_13_nl = MUX_s_1_2_2(or_648_nl, (fsm_output[2]), or_646_nl);
  assign and_641_nl = and_dcpl_72 & and_dcpl_61 & or_dcpl_165;
  assign or_653_nl = (while_if_for_2_for_1_acc_1_tmp[1:0]!=2'b01) | nand_19_cse;
  assign or_651_nl = exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b1101);
  assign mux_15_nl = MUX_s_1_2_2(or_653_nl, (fsm_output[2]), or_651_nl);
  assign and_648_nl = and_dcpl_72 & and_dcpl_65 & or_dcpl_165;
  assign or_656_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b1110);
  assign nor_94_nl = ~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b1110));
  assign mux_17_nl = MUX_s_1_2_2((fsm_output[2]), or_656_nl, nor_94_nl);
  assign and_655_nl = and_dcpl_63 & and_dcpl_65 & or_dcpl_165;
  assign or_659_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b0010);
  assign nor_96_nl = ~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b0010));
  assign mux_19_nl = MUX_s_1_2_2((fsm_output[2]), or_659_nl, nor_96_nl);
  assign and_662_nl = and_dcpl_63 & and_dcpl_69 & or_dcpl_165;
  assign or_662_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b0011);
  assign nor_97_nl = ~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b0011));
  assign mux_21_nl = MUX_s_1_2_2((fsm_output[2]), or_662_nl, nor_97_nl);
  assign and_669_nl = and_dcpl_78 & and_dcpl_71 & or_dcpl_165;
  assign or_666_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b0100);
  assign or_665_nl = exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b0100);
  assign mux_23_nl = MUX_s_1_2_2(or_666_nl, (fsm_output[2]), or_665_nl);
  assign and_676_nl = and_dcpl_78 & and_dcpl_61 & or_dcpl_165;
  assign or_670_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b0101);
  assign or_669_nl = exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b0101);
  assign mux_25_nl = MUX_s_1_2_2(or_670_nl, (fsm_output[2]), or_669_nl);
  assign and_683_nl = and_dcpl_78 & and_dcpl_65 & or_dcpl_165;
  assign or_673_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b0110);
  assign nor_98_nl = ~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b0110));
  assign mux_27_nl = MUX_s_1_2_2((fsm_output[2]), or_673_nl, nor_98_nl);
  assign and_690_nl = and_dcpl_78 & and_dcpl_69 & or_dcpl_165;
  assign nand_22_nl = ~((while_if_for_2_for_1_acc_1_tmp==4'b0111));
  assign nor_99_nl = ~(exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b0111));
  assign mux_29_nl = MUX_s_1_2_2((fsm_output[2]), nand_22_nl, nor_99_nl);
  assign and_697_nl = and_dcpl_67 & and_dcpl_71 & or_dcpl_165;
  assign or_681_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b1000);
  assign or_679_nl = exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b1000);
  assign mux_31_nl = MUX_s_1_2_2(or_681_nl, (fsm_output[2]), or_679_nl);
  assign and_704_nl = and_dcpl_67 & and_dcpl_61 & or_dcpl_165;
  assign or_686_nl = (while_if_for_2_for_1_acc_1_tmp!=4'b1001);
  assign or_684_nl = exit_while_if_for_1_for_1_sva | (while_if_for_1_for_1_n_3_0_sva!=4'b1001);
  assign mux_33_nl = MUX_s_1_2_2(or_686_nl, (fsm_output[2]), or_684_nl);
  assign and_711_nl = in_equal_1_cse & (fsm_output[7]);
  assign and_718_nl = in_equal_2_cse & (fsm_output[7]);
  assign and_725_nl = in_equal_3_cse & (fsm_output[7]);
  assign in_or_14_nl = (and_dcpl_63 & and_dcpl_71 & (out_or_cse | (fsm_output[16])))
      | (fsm_output[21]);
  assign while_if_for_4_not_3_nl = ~ while_if_for_4_and_tmp_1_sva_mx0w0;
  assign while_if_for_4_and_4_nl = MUX_v_16_2_2(16'b0000000000000000, out_10_lpi_2,
      while_if_for_4_not_3_nl);
  assign or_534_nl = (in_equal_2_cse & (fsm_output[17])) | and_753_cse;
  assign while_if_for_4_not_4_nl = ~ while_if_for_4_and_tmp_sva_mx0w0;
  assign while_if_for_4_and_5_nl = MUX_v_16_2_2(16'b0000000000000000, out_11_lpi_2,
      while_if_for_4_not_4_nl);
  assign or_543_nl = (in_equal_3_cse & (fsm_output[17])) | and_774_cse;
  assign while_if_for_for_b_while_if_for_for_b_mux_nl = MUX_v_2_2_2((z_out[1:0]),
      (while_if_for_4_acc_1_cse_1_sva[1:0]), fsm_output[23]);
  assign nor_62_nl = ~((fsm_output[2]) | (fsm_output[9]) | (fsm_output[14]) | (fsm_output[19])
      | ((z_out[2]) & (fsm_output[4])));
  assign regwr_data_not_nl = ~ regwr_data_1_sva_mx0c0;
  assign and_806_nl = in_equal_cse & or_dcpl_204;
  assign or_558_nl = (in_equal_cse & (fsm_output[17])) | and_809_cse;
  assign mux1h_nl = MUX1HOT_v_16_3_2(out_1_lpi_2, while_if_for_3_for_while_if_for_3_for_acc_1_ctmp_sva,
      out_12_sva, {and_806_nl , or_558_nl , (fsm_output[19])});
  assign nor_61_nl = ~((~((~(or_dcpl_55 | (fsm_output[15]))) | while_if_for_1_while_if_for_1_or_1_cse))
      | ((z_out[2]) & (fsm_output[20])));
  assign or_718_nl = (fsm_output[17]) | (fsm_output[12]) | (fsm_output[7]);
  assign mux_37_nl = MUX_s_1_2_2(mux_tmp_36, or_tmp_432, or_718_nl);
  assign mux_38_nl = MUX_s_1_2_2(mux_37_nl, mux_tmp_36, while_if_for_1_while_if_for_1_or_1_cse);
  assign mux_39_nl = MUX_s_1_2_2((~ mux_38_nl), or_tmp_433, or_716_cse);
  assign mux_35_nl = MUX_s_1_2_2((~ or_tmp_432), or_tmp_433, or_716_cse);
  assign mux_40_nl = MUX_s_1_2_2(mux_39_nl, mux_35_nl, fsm_output[19]);
  assign while_if_for_2_for_nor_nl = ~(MUX_v_4_2_2(while_if_for_2_for_1_acc_1_tmp,
      4'b1111, exit_while_if_for_1_for_1_sva));
  assign in_and_nl = in_equal_cse & (fsm_output[5]);
  assign in_and_1_nl = in_equal_1_cse & (fsm_output[5]);
  assign in_and_2_nl = in_equal_2_cse & (fsm_output[5]);
  assign in_and_3_nl = in_equal_3_cse & (fsm_output[5]);
  assign in_and_4_nl = in_equal_cse & (fsm_output[10]);
  assign in_and_5_nl = in_equal_1_cse & (fsm_output[10]);
  assign in_and_6_nl = in_equal_2_cse & (fsm_output[10]);
  assign in_and_7_nl = in_equal_3_cse & (fsm_output[10]);
  assign in_and_8_nl = in_equal_cse & (fsm_output[15]);
  assign in_and_9_nl = in_equal_1_cse & (fsm_output[15]);
  assign in_and_10_nl = in_equal_2_cse & (fsm_output[15]);
  assign in_and_11_nl = in_equal_3_cse & (fsm_output[15]);
  assign in_and_12_nl = in_equal_cse & (fsm_output[20]);
  assign in_and_13_nl = in_equal_1_cse & (fsm_output[20]);
  assign in_and_14_nl = in_equal_2_cse & (fsm_output[20]);
  assign in_and_15_nl = in_equal_3_cse & (fsm_output[20]);
  assign and_846_nl = in_equal_1_cse & (fsm_output[12]);
  assign and_853_nl = in_equal_2_cse & (fsm_output[12]);
  assign and_860_nl = in_equal_3_cse & (fsm_output[12]);
  assign while_if_for_1_for_nor_1_nl = ~((fsm_output[3]) | or_601_ssc | (fsm_output[20]));
  assign while_if_for_1_for_while_if_for_1_for_and_1_nl = MUX_v_2_2_2(2'b00, (while_if_for_1_for_m_4_0_sva_1_3_0[3:2]),
      while_if_for_1_for_nor_1_nl);
  assign while_if_for_1_for_or_1_nl = or_601_ssc | (fsm_output[20]);
  assign while_if_for_1_for_mux1h_1_nl = MUX1HOT_v_2_3_2((while_if_for_1_for_m_4_0_sva_1_3_0[1:0]),
      while_if_for_for_b_2_0_sva_1_0, while_if_for_1_j_2_0_sva_1_0, {or_633_cse ,
      (fsm_output[3]) , while_if_for_1_for_or_1_nl});
  assign nl_z_out = conv_u2u_4_5({while_if_for_1_for_while_if_for_1_for_and_1_nl
      , while_if_for_1_for_mux1h_1_nl}) + 5'b00001;
  assign z_out = nl_z_out[4:0];
  assign or_719_nl = (fsm_output[16]) | (fsm_output[18]);
  assign while_if_for_4_for_mux_39_nl = MUX_v_2_2_2((while_if_for_4_acc_1_cse_1_sva[1:0]),
      while_if_for_1_j_2_0_sva_1_0, or_719_nl);
  assign z_out_4 = MUX_v_16_4_2(out_0_lpi_2, out_1_lpi_2, out_10_lpi_2, out_11_lpi_2,
      while_if_for_4_for_mux_39_nl);

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_16_2;
    input [15:0] input_15;
    input [15:0] input_14;
    input [15:0] input_13;
    input [15:0] input_12;
    input [15:0] input_11;
    input [15:0] input_10;
    input [15:0] input_9;
    input [15:0] input_8;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [15:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    result = result | (input_8 & {16{sel[8]}});
    result = result | (input_9 & {16{sel[9]}});
    result = result | (input_10 & {16{sel[10]}});
    result = result | (input_11 & {16{sel[11]}});
    result = result | (input_12 & {16{sel[12]}});
    result = result | (input_13 & {16{sel[13]}});
    result = result | (input_14 & {16{sel[14]}});
    result = result | (input_15 & {16{sel[15]}});
    MUX1HOT_v_16_16_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_8_2;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [7:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    MUX1HOT_v_16_8_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_9_2;
    input [15:0] input_8;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [8:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    result = result | (input_8 & {16{sel[8]}});
    MUX1HOT_v_16_9_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_16_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_16_16_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_16_2x0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_16_16_2x0 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_4_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [1:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_16_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi (
  clk, reset_bar, if_axi_wr_b_val, if_axi_wr_b_rdy, if_axi_wr_b_msg, run_wen, run_wten,
      if_axi_wr_b_Push_mioi_oswt_unreg, if_axi_wr_b_Push_mioi_bawt, if_axi_wr_b_Push_mioi_iswt0,
      if_axi_wr_b_Push_mioi_wen_comp, if_axi_wr_b_Push_mioi_idat
);
  input clk;
  input reset_bar;
  output if_axi_wr_b_val;
  input if_axi_wr_b_rdy;
  output [5:0] if_axi_wr_b_msg;
  input run_wen;
  input run_wten;
  input if_axi_wr_b_Push_mioi_oswt_unreg;
  output if_axi_wr_b_Push_mioi_bawt;
  input if_axi_wr_b_Push_mioi_iswt0;
  output if_axi_wr_b_Push_mioi_wen_comp;
  input [5:0] if_axi_wr_b_Push_mioi_idat;


  // Interconnect Declarations
  wire if_axi_wr_b_Push_mioi_biwt;
  wire if_axi_wr_b_Push_mioi_bdwt;
  wire if_axi_wr_b_Push_mioi_ivld_run_sct;
  wire if_axi_wr_b_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  wire [5:0] nl_if_axi_wr_b_Push_mioi_idat;
  assign nl_if_axi_wr_b_Push_mioi_idat = {(if_axi_wr_b_Push_mioi_idat[5]) , 1'b0
      , (if_axi_wr_b_Push_mioi_idat[3:0])};
  ccs_out_wait_v1 #(.rscid(32'sd26),
  .width(32'sd6)) if_axi_wr_b_Push_mioi (
      .vld(if_axi_wr_b_val),
      .rdy(if_axi_wr_b_rdy),
      .dat(if_axi_wr_b_msg),
      .ivld(if_axi_wr_b_Push_mioi_ivld_run_sct),
      .irdy(if_axi_wr_b_Push_mioi_irdy),
      .idat(nl_if_axi_wr_b_Push_mioi_idat[5:0])
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_if_axi_wr_b_Push_mio_wait_ctrl
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_if_axi_wr_b_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_wr_b_Push_mioi_oswt_unreg(if_axi_wr_b_Push_mioi_oswt_unreg),
      .if_axi_wr_b_Push_mioi_iswt0(if_axi_wr_b_Push_mioi_iswt0),
      .if_axi_wr_b_Push_mioi_biwt(if_axi_wr_b_Push_mioi_biwt),
      .if_axi_wr_b_Push_mioi_bdwt(if_axi_wr_b_Push_mioi_bdwt),
      .if_axi_wr_b_Push_mioi_ivld_run_sct(if_axi_wr_b_Push_mioi_ivld_run_sct),
      .if_axi_wr_b_Push_mioi_irdy(if_axi_wr_b_Push_mioi_irdy)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_if_axi_wr_b_Push_mio_wait_dp
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_if_axi_wr_b_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_wr_b_Push_mioi_oswt_unreg(if_axi_wr_b_Push_mioi_oswt_unreg),
      .if_axi_wr_b_Push_mioi_bawt(if_axi_wr_b_Push_mioi_bawt),
      .if_axi_wr_b_Push_mioi_wen_comp(if_axi_wr_b_Push_mioi_wen_comp),
      .if_axi_wr_b_Push_mioi_biwt(if_axi_wr_b_Push_mioi_biwt),
      .if_axi_wr_b_Push_mioi_bdwt(if_axi_wr_b_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi (
  clk, reset_bar, if_axi_wr_w_val, if_axi_wr_w_rdy, if_axi_wr_w_msg, run_wen, run_wten,
      if_axi_wr_w_PopNB_mioi_oswt_unreg, if_axi_wr_w_PopNB_mioi_bawt, if_axi_wr_w_PopNB_mioi_iswt0,
      if_axi_wr_w_PopNB_mioi_ivld_mxwt, if_axi_wr_w_PopNB_mioi_idat_mxwt
);
  input clk;
  input reset_bar;
  input if_axi_wr_w_val;
  output if_axi_wr_w_rdy;
  input [72:0] if_axi_wr_w_msg;
  input run_wen;
  input run_wten;
  input if_axi_wr_w_PopNB_mioi_oswt_unreg;
  output if_axi_wr_w_PopNB_mioi_bawt;
  input if_axi_wr_w_PopNB_mioi_iswt0;
  output if_axi_wr_w_PopNB_mioi_ivld_mxwt;
  output [72:0] if_axi_wr_w_PopNB_mioi_idat_mxwt;


  // Interconnect Declarations
  wire if_axi_wr_w_PopNB_mioi_biwt;
  wire if_axi_wr_w_PopNB_mioi_bdwt;
  wire if_axi_wr_w_PopNB_mioi_ivld;
  wire [72:0] if_axi_wr_w_PopNB_mioi_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd25),
  .width(32'sd73)) if_axi_wr_w_PopNB_mioi (
      .vld(if_axi_wr_w_val),
      .rdy(if_axi_wr_w_rdy),
      .dat(if_axi_wr_w_msg),
      .ivld(if_axi_wr_w_PopNB_mioi_ivld),
      .irdy(if_axi_wr_w_PopNB_mioi_biwt),
      .idat(if_axi_wr_w_PopNB_mioi_idat)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_if_axi_wr_w_PopNB_mio_wait_ctrl
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_if_axi_wr_w_PopNB_mio_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_wr_w_PopNB_mioi_oswt_unreg(if_axi_wr_w_PopNB_mioi_oswt_unreg),
      .if_axi_wr_w_PopNB_mioi_iswt0(if_axi_wr_w_PopNB_mioi_iswt0),
      .if_axi_wr_w_PopNB_mioi_biwt(if_axi_wr_w_PopNB_mioi_biwt),
      .if_axi_wr_w_PopNB_mioi_bdwt(if_axi_wr_w_PopNB_mioi_bdwt)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_if_axi_wr_w_PopNB_mio_wait_dp
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_if_axi_wr_w_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_wr_w_PopNB_mioi_bawt(if_axi_wr_w_PopNB_mioi_bawt),
      .if_axi_wr_w_PopNB_mioi_ivld_mxwt(if_axi_wr_w_PopNB_mioi_ivld_mxwt),
      .if_axi_wr_w_PopNB_mioi_idat_mxwt(if_axi_wr_w_PopNB_mioi_idat_mxwt),
      .if_axi_wr_w_PopNB_mioi_biwt(if_axi_wr_w_PopNB_mioi_biwt),
      .if_axi_wr_w_PopNB_mioi_bdwt(if_axi_wr_w_PopNB_mioi_bdwt),
      .if_axi_wr_w_PopNB_mioi_ivld(if_axi_wr_w_PopNB_mioi_ivld),
      .if_axi_wr_w_PopNB_mioi_idat(if_axi_wr_w_PopNB_mioi_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi (
  clk, reset_bar, if_axi_rd_r_val, if_axi_rd_r_rdy, if_axi_rd_r_msg, run_wen, run_wten,
      if_axi_rd_r_Push_mioi_oswt_unreg, if_axi_rd_r_Push_mioi_bawt, if_axi_rd_r_Push_mioi_iswt0,
      if_axi_rd_r_Push_mioi_wen_comp, if_axi_rd_r_Push_mioi_idat
);
  input clk;
  input reset_bar;
  output if_axi_rd_r_val;
  input if_axi_rd_r_rdy;
  output [70:0] if_axi_rd_r_msg;
  input run_wen;
  input run_wten;
  input if_axi_rd_r_Push_mioi_oswt_unreg;
  output if_axi_rd_r_Push_mioi_bawt;
  input if_axi_rd_r_Push_mioi_iswt0;
  output if_axi_rd_r_Push_mioi_wen_comp;
  input [70:0] if_axi_rd_r_Push_mioi_idat;


  // Interconnect Declarations
  wire if_axi_rd_r_Push_mioi_biwt;
  wire if_axi_rd_r_Push_mioi_bdwt;
  wire if_axi_rd_r_Push_mioi_ivld_run_sct;
  wire if_axi_rd_r_Push_mioi_irdy;


  // Interconnect Declarations for Component Instantiations 
  wire [70:0] nl_if_axi_rd_r_Push_mioi_idat;
  assign nl_if_axi_rd_r_Push_mioi_idat = {(if_axi_rd_r_Push_mioi_idat[70:69]) , 1'b0
      , (if_axi_rd_r_Push_mioi_idat[67:0])};
  ccs_out_wait_v1 #(.rscid(32'sd24),
  .width(32'sd71)) if_axi_rd_r_Push_mioi (
      .vld(if_axi_rd_r_val),
      .rdy(if_axi_rd_r_rdy),
      .dat(if_axi_rd_r_msg),
      .ivld(if_axi_rd_r_Push_mioi_ivld_run_sct),
      .irdy(if_axi_rd_r_Push_mioi_irdy),
      .idat(nl_if_axi_rd_r_Push_mioi_idat[70:0])
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_if_axi_rd_r_Push_mio_wait_ctrl
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_if_axi_rd_r_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_rd_r_Push_mioi_oswt_unreg(if_axi_rd_r_Push_mioi_oswt_unreg),
      .if_axi_rd_r_Push_mioi_iswt0(if_axi_rd_r_Push_mioi_iswt0),
      .if_axi_rd_r_Push_mioi_biwt(if_axi_rd_r_Push_mioi_biwt),
      .if_axi_rd_r_Push_mioi_bdwt(if_axi_rd_r_Push_mioi_bdwt),
      .if_axi_rd_r_Push_mioi_ivld_run_sct(if_axi_rd_r_Push_mioi_ivld_run_sct),
      .if_axi_rd_r_Push_mioi_irdy(if_axi_rd_r_Push_mioi_irdy)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_if_axi_rd_r_Push_mio_wait_dp
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_if_axi_rd_r_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_rd_r_Push_mioi_oswt_unreg(if_axi_rd_r_Push_mioi_oswt_unreg),
      .if_axi_rd_r_Push_mioi_bawt(if_axi_rd_r_Push_mioi_bawt),
      .if_axi_rd_r_Push_mioi_wen_comp(if_axi_rd_r_Push_mioi_wen_comp),
      .if_axi_rd_r_Push_mioi_biwt(if_axi_rd_r_Push_mioi_biwt),
      .if_axi_rd_r_Push_mioi_bdwt(if_axi_rd_r_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi (
  clk, reset_bar, regIn_val, regIn_rdy, regIn_msg, run_wen, run_wten, regIn_PopNB_mioi_oswt_unreg,
      regIn_PopNB_mioi_bawt, regIn_PopNB_mioi_iswt0, regIn_PopNB_mioi_ivld_mxwt,
      regIn_PopNB_mioi_idat_mxwt
);
  input clk;
  input reset_bar;
  input regIn_val;
  output regIn_rdy;
  input [70:0] regIn_msg;
  input run_wen;
  input run_wten;
  input regIn_PopNB_mioi_oswt_unreg;
  output regIn_PopNB_mioi_bawt;
  input regIn_PopNB_mioi_iswt0;
  output regIn_PopNB_mioi_ivld_mxwt;
  output [67:0] regIn_PopNB_mioi_idat_mxwt;


  // Interconnect Declarations
  wire regIn_PopNB_mioi_biwt;
  wire regIn_PopNB_mioi_bdwt;
  wire regIn_PopNB_mioi_ivld;
  wire [70:0] regIn_PopNB_mioi_idat;
  wire [67:0] regIn_PopNB_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd23),
  .width(32'sd71)) regIn_PopNB_mioi (
      .vld(regIn_val),
      .rdy(regIn_rdy),
      .dat(regIn_msg),
      .ivld(regIn_PopNB_mioi_ivld),
      .irdy(regIn_PopNB_mioi_biwt),
      .idat(regIn_PopNB_mioi_idat)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_regIn_PopNB_mio_wait_ctrl
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_regIn_PopNB_mio_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .regIn_PopNB_mioi_oswt_unreg(regIn_PopNB_mioi_oswt_unreg),
      .regIn_PopNB_mioi_iswt0(regIn_PopNB_mioi_iswt0),
      .regIn_PopNB_mioi_biwt(regIn_PopNB_mioi_biwt),
      .regIn_PopNB_mioi_bdwt(regIn_PopNB_mioi_bdwt)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_regIn_PopNB_mio_wait_dp
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_regIn_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .regIn_PopNB_mioi_bawt(regIn_PopNB_mioi_bawt),
      .regIn_PopNB_mioi_ivld_mxwt(regIn_PopNB_mioi_ivld_mxwt),
      .regIn_PopNB_mioi_idat_mxwt(regIn_PopNB_mioi_idat_mxwt_pconst),
      .regIn_PopNB_mioi_biwt(regIn_PopNB_mioi_biwt),
      .regIn_PopNB_mioi_bdwt(regIn_PopNB_mioi_bdwt),
      .regIn_PopNB_mioi_ivld(regIn_PopNB_mioi_ivld),
      .regIn_PopNB_mioi_idat(regIn_PopNB_mioi_idat)
    );
  assign regIn_PopNB_mioi_idat_mxwt = regIn_PopNB_mioi_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi (
  clk, reset_bar, if_axi_wr_aw_val, if_axi_wr_aw_rdy, if_axi_wr_aw_msg, run_wen,
      run_wten, if_axi_wr_aw_PopNB_mioi_oswt_unreg, if_axi_wr_aw_PopNB_mioi_bawt,
      if_axi_wr_aw_PopNB_mioi_iswt0, if_axi_wr_aw_PopNB_mioi_ivld_mxwt, if_axi_wr_aw_PopNB_mioi_idat_mxwt
);
  input clk;
  input reset_bar;
  input if_axi_wr_aw_val;
  output if_axi_wr_aw_rdy;
  input [43:0] if_axi_wr_aw_msg;
  input run_wen;
  input run_wten;
  input if_axi_wr_aw_PopNB_mioi_oswt_unreg;
  output if_axi_wr_aw_PopNB_mioi_bawt;
  input if_axi_wr_aw_PopNB_mioi_iswt0;
  output if_axi_wr_aw_PopNB_mioi_ivld_mxwt;
  output [19:0] if_axi_wr_aw_PopNB_mioi_idat_mxwt;


  // Interconnect Declarations
  wire if_axi_wr_aw_PopNB_mioi_biwt;
  wire if_axi_wr_aw_PopNB_mioi_bdwt;
  wire if_axi_wr_aw_PopNB_mioi_ivld;
  wire [43:0] if_axi_wr_aw_PopNB_mioi_idat;
  wire [19:0] if_axi_wr_aw_PopNB_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd22),
  .width(32'sd44)) if_axi_wr_aw_PopNB_mioi (
      .vld(if_axi_wr_aw_val),
      .rdy(if_axi_wr_aw_rdy),
      .dat(if_axi_wr_aw_msg),
      .ivld(if_axi_wr_aw_PopNB_mioi_ivld),
      .irdy(if_axi_wr_aw_PopNB_mioi_biwt),
      .idat(if_axi_wr_aw_PopNB_mioi_idat)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_if_axi_wr_aw_PopNB_mio_wait_ctrl
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_if_axi_wr_aw_PopNB_mio_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_wr_aw_PopNB_mioi_oswt_unreg(if_axi_wr_aw_PopNB_mioi_oswt_unreg),
      .if_axi_wr_aw_PopNB_mioi_iswt0(if_axi_wr_aw_PopNB_mioi_iswt0),
      .if_axi_wr_aw_PopNB_mioi_biwt(if_axi_wr_aw_PopNB_mioi_biwt),
      .if_axi_wr_aw_PopNB_mioi_bdwt(if_axi_wr_aw_PopNB_mioi_bdwt)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_if_axi_wr_aw_PopNB_mio_wait_dp
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_if_axi_wr_aw_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_wr_aw_PopNB_mioi_bawt(if_axi_wr_aw_PopNB_mioi_bawt),
      .if_axi_wr_aw_PopNB_mioi_ivld_mxwt(if_axi_wr_aw_PopNB_mioi_ivld_mxwt),
      .if_axi_wr_aw_PopNB_mioi_idat_mxwt(if_axi_wr_aw_PopNB_mioi_idat_mxwt_pconst),
      .if_axi_wr_aw_PopNB_mioi_biwt(if_axi_wr_aw_PopNB_mioi_biwt),
      .if_axi_wr_aw_PopNB_mioi_bdwt(if_axi_wr_aw_PopNB_mioi_bdwt),
      .if_axi_wr_aw_PopNB_mioi_ivld(if_axi_wr_aw_PopNB_mioi_ivld),
      .if_axi_wr_aw_PopNB_mioi_idat(if_axi_wr_aw_PopNB_mioi_idat)
    );
  assign if_axi_wr_aw_PopNB_mioi_idat_mxwt = if_axi_wr_aw_PopNB_mioi_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi (
  clk, reset_bar, if_axi_rd_ar_val, if_axi_rd_ar_rdy, if_axi_rd_ar_msg, run_wen,
      run_wten, if_axi_rd_ar_PopNB_mioi_oswt_unreg, if_axi_rd_ar_PopNB_mioi_bawt,
      if_axi_rd_ar_PopNB_mioi_iswt0, if_axi_rd_ar_PopNB_mioi_ivld_mxwt, if_axi_rd_ar_PopNB_mioi_idat_mxwt
);
  input clk;
  input reset_bar;
  input if_axi_rd_ar_val;
  output if_axi_rd_ar_rdy;
  input [43:0] if_axi_rd_ar_msg;
  input run_wen;
  input run_wten;
  input if_axi_rd_ar_PopNB_mioi_oswt_unreg;
  output if_axi_rd_ar_PopNB_mioi_bawt;
  input if_axi_rd_ar_PopNB_mioi_iswt0;
  output if_axi_rd_ar_PopNB_mioi_ivld_mxwt;
  output [27:0] if_axi_rd_ar_PopNB_mioi_idat_mxwt;


  // Interconnect Declarations
  wire if_axi_rd_ar_PopNB_mioi_biwt;
  wire if_axi_rd_ar_PopNB_mioi_bdwt;
  wire if_axi_rd_ar_PopNB_mioi_ivld;
  wire [43:0] if_axi_rd_ar_PopNB_mioi_idat;
  wire [27:0] if_axi_rd_ar_PopNB_mioi_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd21),
  .width(32'sd44)) if_axi_rd_ar_PopNB_mioi (
      .vld(if_axi_rd_ar_val),
      .rdy(if_axi_rd_ar_rdy),
      .dat(if_axi_rd_ar_msg),
      .ivld(if_axi_rd_ar_PopNB_mioi_ivld),
      .irdy(if_axi_rd_ar_PopNB_mioi_biwt),
      .idat(if_axi_rd_ar_PopNB_mioi_idat)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_if_axi_rd_ar_PopNB_mio_wait_ctrl
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_if_axi_rd_ar_PopNB_mio_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_rd_ar_PopNB_mioi_oswt_unreg(if_axi_rd_ar_PopNB_mioi_oswt_unreg),
      .if_axi_rd_ar_PopNB_mioi_iswt0(if_axi_rd_ar_PopNB_mioi_iswt0),
      .if_axi_rd_ar_PopNB_mioi_biwt(if_axi_rd_ar_PopNB_mioi_biwt),
      .if_axi_rd_ar_PopNB_mioi_bdwt(if_axi_rd_ar_PopNB_mioi_bdwt)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_if_axi_rd_ar_PopNB_mio_wait_dp
      AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_if_axi_rd_ar_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_rd_ar_PopNB_mioi_bawt(if_axi_rd_ar_PopNB_mioi_bawt),
      .if_axi_rd_ar_PopNB_mioi_ivld_mxwt(if_axi_rd_ar_PopNB_mioi_ivld_mxwt),
      .if_axi_rd_ar_PopNB_mioi_idat_mxwt(if_axi_rd_ar_PopNB_mioi_idat_mxwt_pconst),
      .if_axi_rd_ar_PopNB_mioi_biwt(if_axi_rd_ar_PopNB_mioi_biwt),
      .if_axi_rd_ar_PopNB_mioi_bdwt(if_axi_rd_ar_PopNB_mioi_bdwt),
      .if_axi_rd_ar_PopNB_mioi_ivld(if_axi_rd_ar_PopNB_mioi_ivld),
      .if_axi_rd_ar_PopNB_mioi_idat(if_axi_rd_ar_PopNB_mioi_idat)
    );
  assign if_axi_rd_ar_PopNB_mioi_idat_mxwt = if_axi_rd_ar_PopNB_mioi_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Accelerator_run
// ------------------------------------------------------------------


module Accelerator_run (
  clk, reset_bar, regOut_chan_0, regOut_chan_1, regOut_chan_2, regOut_chan_3, regOut_chan_4,
      regOut_chan_5, regOut_chan_6, regOut_chan_7, regOut_chan_8, regOut_chan_9,
      regIn_chan_val, regIn_chan_rdy, regIn_chan_msg
);
  input clk;
  input reset_bar;
  input [63:0] regOut_chan_0;
  input [63:0] regOut_chan_1;
  input [63:0] regOut_chan_2;
  input [63:0] regOut_chan_3;
  input [63:0] regOut_chan_4;
  input [63:0] regOut_chan_5;
  input [63:0] regOut_chan_6;
  input [63:0] regOut_chan_7;
  input [63:0] regOut_chan_8;
  input [63:0] regOut_chan_9;
  output regIn_chan_val;
  input regIn_chan_rdy;
  output [70:0] regIn_chan_msg;


  // Interconnect Declarations
  wire regIn_chan_PushNB_mioi_ivld;
  wire regIn_chan_PushNB_mioi_irdy;
  wire [70:0] regIn_chan_PushNB_mioi_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd35),
  .width(32'sd71)) regIn_chan_PushNB_mioi (
      .vld(regIn_chan_val),
      .rdy(regIn_chan_rdy),
      .dat(regIn_chan_msg),
      .ivld(regIn_chan_PushNB_mioi_ivld),
      .irdy(regIn_chan_PushNB_mioi_irdy),
      .idat(regIn_chan_PushNB_mioi_idat)
    );
  Accelerator_run_run Accelerator_run_run_inst (
      .clk(clk),
      .reset_bar(reset_bar),
      .regOut_chan_1(regOut_chan_1),
      .regOut_chan_2(regOut_chan_2),
      .regOut_chan_3(regOut_chan_3),
      .regOut_chan_4(regOut_chan_4),
      .regOut_chan_5(regOut_chan_5),
      .regOut_chan_6(regOut_chan_6),
      .regOut_chan_7(regOut_chan_7),
      .regOut_chan_8(regOut_chan_8),
      .regOut_chan_9(regOut_chan_9),
      .regIn_chan_PushNB_mioi_ivld(regIn_chan_PushNB_mioi_ivld),
      .regIn_chan_PushNB_mioi_irdy(regIn_chan_PushNB_mioi_irdy),
      .regIn_chan_PushNB_mioi_idat(regIn_chan_PushNB_mioi_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16_run
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16_run (
  clk, reset_bar, if_axi_rd_ar_val, if_axi_rd_ar_rdy, if_axi_rd_ar_msg, if_axi_rd_r_val,
      if_axi_rd_r_rdy, if_axi_rd_r_msg, if_axi_wr_aw_val, if_axi_wr_aw_rdy, if_axi_wr_aw_msg,
      if_axi_wr_w_val, if_axi_wr_w_rdy, if_axi_wr_w_msg, if_axi_wr_b_val, if_axi_wr_b_rdy,
      if_axi_wr_b_msg, baseAddr, regOut_0, regOut_1, regOut_2, regOut_3, regOut_4,
      regOut_5, regOut_6, regOut_7, regOut_8, regOut_9, regOut_10, regOut_11, regOut_12,
      regOut_13, regIn_val, regIn_rdy, regIn_msg
);
  input clk;
  input reset_bar;
  input if_axi_rd_ar_val;
  output if_axi_rd_ar_rdy;
  input [43:0] if_axi_rd_ar_msg;
  output if_axi_rd_r_val;
  input if_axi_rd_r_rdy;
  output [70:0] if_axi_rd_r_msg;
  input if_axi_wr_aw_val;
  output if_axi_wr_aw_rdy;
  input [43:0] if_axi_wr_aw_msg;
  input if_axi_wr_w_val;
  output if_axi_wr_w_rdy;
  input [72:0] if_axi_wr_w_msg;
  output if_axi_wr_b_val;
  input if_axi_wr_b_rdy;
  output [5:0] if_axi_wr_b_msg;
  input [15:0] baseAddr;
  output [63:0] regOut_0;
  reg [63:0] regOut_0;
  output [63:0] regOut_1;
  reg [63:0] regOut_1;
  output [63:0] regOut_2;
  reg [63:0] regOut_2;
  output [63:0] regOut_3;
  reg [63:0] regOut_3;
  output [63:0] regOut_4;
  output [63:0] regOut_5;
  reg [63:0] regOut_5;
  output [63:0] regOut_6;
  reg [63:0] regOut_6;
  output [63:0] regOut_7;
  reg [63:0] regOut_7;
  output [63:0] regOut_8;
  output [63:0] regOut_9;
  reg [63:0] regOut_9;
  output [63:0] regOut_10;
  reg [63:0] regOut_10;
  output [63:0] regOut_11;
  reg [63:0] regOut_11;
  output [63:0] regOut_12;
  reg [63:0] regOut_12;
  output [63:0] regOut_13;
  reg [63:0] regOut_13;
  input regIn_val;
  output regIn_rdy;
  input [70:0] regIn_msg;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire if_axi_rd_ar_PopNB_mioi_bawt;
  reg if_axi_rd_ar_PopNB_mioi_iswt0;
  wire if_axi_rd_ar_PopNB_mioi_ivld_mxwt;
  wire [27:0] if_axi_rd_ar_PopNB_mioi_idat_mxwt;
  wire if_axi_wr_aw_PopNB_mioi_bawt;
  reg if_axi_wr_aw_PopNB_mioi_iswt0;
  wire if_axi_wr_aw_PopNB_mioi_ivld_mxwt;
  wire [19:0] if_axi_wr_aw_PopNB_mioi_idat_mxwt;
  wire regIn_PopNB_mioi_bawt;
  reg regIn_PopNB_mioi_iswt0;
  wire regIn_PopNB_mioi_ivld_mxwt;
  wire [67:0] regIn_PopNB_mioi_idat_mxwt;
  wire if_axi_rd_r_Push_mioi_bawt;
  reg if_axi_rd_r_Push_mioi_iswt0;
  wire if_axi_rd_r_Push_mioi_wen_comp;
  wire if_axi_wr_w_PopNB_mioi_bawt;
  reg if_axi_wr_w_PopNB_mioi_iswt0;
  wire if_axi_wr_w_PopNB_mioi_ivld_mxwt;
  wire [72:0] if_axi_wr_w_PopNB_mioi_idat_mxwt;
  wire if_axi_wr_b_Push_mioi_bawt;
  reg if_axi_wr_b_Push_mioi_iswt0;
  wire if_axi_wr_b_Push_mioi_wen_comp;
  reg if_axi_rd_r_Push_mioi_idat_70;
  reg if_axi_rd_r_Push_mioi_idat_69;
  reg [63:0] if_axi_rd_r_Push_mioi_idat_67_4;
  reg [3:0] if_axi_rd_r_Push_mioi_idat_3_0;
  reg if_axi_wr_b_Push_mioi_idat_5;
  reg [3:0] if_axi_wr_b_Push_mioi_idat_3_0;
  wire [1:0] fsm_output;
  wire while_while_or_2_tmp;
  wire while_while_or_1_tmp;
  wire while_while_or_tmp;
  wire [7:0] while_mux_17_tmp;
  wire [3:0] while_mux_32_tmp;
  wire and_dcpl;
  wire or_dcpl_2;
  wire or_dcpl_3;
  wire or_dcpl_4;
  wire or_tmp_54;
  wire nand_tmp_10;
  wire mux_tmp_86;
  wire mux_tmp_87;
  wire nand_tmp_14;
  wire or_tmp_70;
  wire nand_tmp_15;
  wire mux_tmp_112;
  wire nand_tmp_19;
  wire or_tmp_86;
  wire nand_tmp_20;
  wire mux_tmp_136;
  wire mux_tmp_143;
  wire or_tmp_103;
  wire mux_tmp_144;
  wire mux_tmp_149;
  wire or_tmp_114;
  wire nand_tmp_26;
  wire mux_tmp_168;
  wire mux_tmp_169;
  wire nand_tmp_30;
  wire or_tmp_129;
  wire nand_tmp_31;
  wire mux_tmp_194;
  wire mux_tmp_195;
  wire nand_tmp_35;
  wire or_tmp_145;
  wire nand_tmp_36;
  wire mux_tmp_220;
  wire mux_tmp_221;
  wire mux_tmp_234;
  wire or_tmp_172;
  wire nand_tmp_42;
  wire mux_tmp_253;
  wire nand_tmp_46;
  wire or_tmp_188;
  wire nand_tmp_47;
  wire mux_tmp_277;
  wire mux_tmp_278;
  wire nand_tmp_51;
  wire or_tmp_204;
  wire nand_tmp_52;
  wire mux_tmp_303;
  wire mux_tmp_304;
  wire nand_tmp_56;
  wire or_dcpl_17;
  wire or_tmp_221;
  wire or_tmp_228;
  wire or_tmp_234;
  wire and_dcpl_19;
  wire and_dcpl_20;
  wire nor_tmp_25;
  wire mux_tmp_364;
  wire or_dcpl_25;
  wire and_dcpl_24;
  wire and_dcpl_25;
  wire and_dcpl_26;
  wire or_dcpl_28;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire or_dcpl_35;
  wire or_dcpl_36;
  wire or_dcpl_38;
  wire or_dcpl_39;
  wire or_tmp_280;
  wire or_tmp_282;
  wire not_tmp_228;
  wire mux_tmp_370;
  wire and_tmp_19;
  wire or_tmp_285;
  wire or_tmp_287;
  wire mux_tmp_373;
  wire nand_tmp_63;
  wire nand_tmp_66;
  wire mux_tmp_378;
  wire or_tmp_292;
  wire mux_tmp_381;
  wire nor_tmp_28;
  wire nor_tmp_30;
  wire and_dcpl_55;
  wire and_dcpl_58;
  wire nand_tmp_71;
  wire and_tmp_21;
  wire or_tmp_311;
  wire or_tmp_315;
  wire or_tmp_322;
  wire and_tmp_26;
  wire nand_tmp_74;
  wire not_tmp_258;
  wire or_dcpl_43;
  wire mux_tmp_423;
  wire and_tmp_32;
  wire mux_tmp_424;
  wire and_tmp_33;
  wire mux_tmp_427;
  wire or_tmp_349;
  wire nand_tmp_80;
  wire mux_tmp_431;
  wire mux_tmp_437;
  wire nand_tmp_85;
  wire and_tmp_36;
  wire mux_tmp_455;
  wire or_tmp_368;
  wire or_tmp_369;
  wire or_tmp_370;
  wire or_tmp_371;
  wire or_tmp_377;
  wire or_tmp_378;
  wire or_tmp_384;
  wire or_tmp_385;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_83;
  wire and_tmp_39;
  wire and_tmp_40;
  wire or_dcpl_51;
  wire and_dcpl_91;
  wire or_dcpl_52;
  wire or_tmp_435;
  wire mux_tmp_519;
  wire and_tmp_60;
  wire and_tmp_61;
  wire mux_tmp_527;
  wire mux_tmp_530;
  wire mux_tmp_545;
  wire or_tmp_439;
  wire or_tmp_456;
  wire mux_tmp_559;
  wire mux_tmp_562;
  wire mux_tmp_575;
  wire and_dcpl_117;
  wire or_dcpl_64;
  wire nand_tmp_98;
  wire and_tmp_70;
  wire and_tmp_71;
  wire and_tmp_72;
  wire and_tmp_75;
  wire and_tmp_76;
  wire or_tmp_509;
  wire or_tmp_510;
  wire mux_tmp_611;
  wire mux_tmp_614;
  wire or_tmp_514;
  wire and_tmp_78;
  wire nand_tmp_102;
  wire nand_tmp_103;
  wire mux_tmp_622;
  wire mux_tmp_633;
  wire mux_tmp_642;
  wire not_tmp_372;
  wire mux_tmp_653;
  wire not_tmp_373;
  wire mux_tmp_656;
  wire or_tmp_529;
  wire and_dcpl_130;
  wire or_tmp_576;
  wire and_256_cse;
  wire select_mask_2_1_sva_dfm_0_mx0;
  wire select_mask_2_1_sva_dfm_1_mx0;
  wire select_mask_0_sva_dfm_mx0;
  wire operator_5_false_operator_5_false_operator_5_false_or_svs_mx1;
  wire nvhls_set_slc_Arbiter_3U_Roundrobin_Mask_nvhls_nvhls_t_2U_nvuint_t_X_temp_2_1_sva_1_1;
  wire arb_pick_priority_4_sva_mx0w0;
  wire nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm_mx0w0;
  wire nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm_mx0w0;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1;
  wire regIn_arb_req_sva_mx1;
  wire arb_pick_priority_3_sva_1;
  wire read_arb_req_sva_mx1;
  wire write_arb_req_sva_mx1;
  reg arb_next_1_2_sva;
  reg arb_next_1_1_sva;
  wire while_or_16_cse_1;
  wire while_or_17_cse_1;
  wire while_or_18_cse_1;
  wire while_or_19_cse_1;
  wire while_or_cse_1;
  wire while_or_14_cse_1;
  wire [7:0] axiRdLen_sva_dfm_1_mx0;
  reg read_arb_req_sva;
  reg while_stage_v_1;
  reg operator_3_false_2_operator_3_false_2_and_svs_st_1;
  reg operator_3_false_1_operator_3_false_1_and_svs_st_1;
  reg while_asn_34_itm_1;
  reg while_asn_30_itm_1;
  reg while_asn_25_itm_1;
  reg while_else_4_if_if_for_equal_tmp_13_1;
  reg while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  wire while_else_4_else_if_and_stg_2_5_sva_1;
  reg operator_3_false_3_operator_3_false_3_and_svs_2;
  reg while_else_4_if_if_for_equal_tmp_12_1;
  wire while_else_4_else_if_and_stg_2_4_sva_1;
  reg while_else_4_if_if_for_equal_tmp_11_1;
  wire while_else_4_else_if_and_stg_2_3_sva_1;
  reg while_else_4_if_if_for_equal_tmp_10_1;
  wire while_else_4_else_if_and_stg_2_2_sva_1;
  reg while_else_4_if_if_for_equal_tmp_9_1;
  wire while_else_4_else_if_and_stg_2_1_sva_1;
  wire while_else_4_else_if_and_stg_2_0_sva_1;
  reg while_else_4_if_if_for_equal_tmp_7_1;
  wire while_else_4_else_if_and_stg_1_3_sva_1;
  reg while_else_4_if_if_for_equal_tmp_6_1;
  wire while_else_4_else_if_and_stg_1_2_sva_1;
  reg while_else_4_if_if_for_equal_tmp_5_1;
  reg while_else_4_if_if_for_equal_tmp_3_1;
  reg operator_3_false_2_operator_3_false_2_and_svs_2;
  reg operator_3_false_1_operator_3_false_1_and_svs_2;
  reg while_else_4_if_if_for_while_else_4_if_if_for_and_13_itm_1;
  reg while_else_4_if_if_for_while_else_4_if_if_for_and_14_itm_1;
  reg [3:0] operator_17_true_return_1_3_0_sva_1;
  reg while_else_4_if_if_for_nor_6_itm_1;
  reg while_else_4_if_if_for_nor_3_itm_1;
  reg while_else_4_if_if_for_nor_1_itm_1;
  reg while_else_4_if_if_for_nor_itm_1;
  wire while_else_4_else_if_and_stg_1_0_sva_1;
  wire while_else_4_else_if_and_stg_1_1_sva_1;
  reg while_stage_v_2;
  reg while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1;
  reg while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1;
  reg operator_3_false_2_operator_3_false_2_and_svs_st_2;
  reg operator_3_false_1_operator_3_false_1_and_svs_st_2;
  wire arb_pick_return_2_1_lpi_1_dfm_1_1_1;
  wire arb_pick_return_2_1_lpi_1_dfm_1_0_1;
  wire arb_pick_return_0_lpi_1_dfm_2;
  reg operator_3_false_1_operator_3_false_1_and_svs_1;
  reg [3:0] regwr_addr_6_3_sva;
  reg operator_3_false_3_operator_3_false_3_and_svs_1;
  reg operator_3_false_3_operator_3_false_3_and_svs_st_1;
  reg operator_3_false_2_operator_3_false_2_and_svs_1;
  reg write_arb_req_sva;
  reg while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  reg [2:0] if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70;
  reg regIn_arb_req_sva;
  reg arb_needs_update_sva;
  reg operator_8_false_operator_8_false_nor_mdf_sva;
  reg select_mask_2_1_sva_1;
  reg select_mask_2_1_sva_0;
  wire arb_pick_if_1_and_tmp_2_mx0w0;
  reg arb_pick_if_1_and_tmp_2;
  wire operator_3_false_operator_3_false_nor_svs_1;
  reg nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm;
  reg nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm;
  wire arb_pick_priority_4_sva_mx1;
  wire arb_pick_if_1_and_stg_1_0_mx0w0;
  reg arb_pick_if_1_and_stg_1_0;
  wire operator_8_false_operator_8_false_nor_mdf_sva_mx1;
  wire if_axi_wr_bwrite_and_cse;
  wire nor_124_cse;
  wire regOut_13_and_cse;
  wire or_28_cse;
  wire or_26_cse;
  wire and_309_cse;
  wire and_312_cse;
  wire and_314_cse;
  wire nor_97_cse;
  wire or_210_cse;
  wire nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_and_1_cse;
  wire regIn_arb_req_and_cse;
  wire select_mask_and_cse;
  wire arb_needs_update_and_cse;
  wire operator_3_false_3_and_cse;
  wire while_and_98_cse;
  wire operator_3_false_2_and_2_cse;
  wire and_352_cse;
  wire or_310_cse;
  wire or_662_cse;
  wire nor_70_cse;
  wire or_673_cse;
  wire nor_81_cse;
  wire while_nand_2_cse;
  wire and_305_cse;
  wire or_234_cse;
  wire nor_116_cse;
  reg [63:0] reg_regOut_8_cse;
  reg [63:0] reg_regOut_4_cse;
  wire arb_next_and_cse;
  wire mux_5_cse;
  wire mux_151_cse;
  wire nor_132_cse;
  wire or_68_cse;
  wire nor_136_cse;
  wire or_100_cse;
  wire or_668_cse;
  wire or_143_cse;
  wire while_stage_en_1_mx0w1;
  wire mux_374_itm;
  wire mux_404_itm;
  wire mux_481_itm;
  wire mux_488_itm;
  wire mux_489_itm;
  wire mux_555_itm;
  wire mux_610_itm;
  wire [16:0] z_out;
  wire [12:0] z_out_1;
  wire [13:0] nl_z_out_1;
  reg [15:0] operator_33_true_return_15_0_sva;
  reg [63:0] reg_6_sva;
  reg [63:0] reg_7_sva;
  reg [63:0] reg_5_sva;
  reg [63:0] reg_9_sva;
  reg [63:0] reg_3_sva;
  reg [63:0] reg_10_sva;
  reg [63:0] reg_2_sva;
  reg [63:0] reg_11_sva;
  reg [63:0] reg_1_sva;
  reg [63:0] reg_12_sva;
  reg [63:0] reg_0_sva;
  reg [63:0] reg_13_sva;
  reg [3:0] axi_rd_req_id_sva;
  reg [63:0] axi_rd_resp_data_sva;
  reg [3:0] axi_wr_req_addr_id_sva;
  reg [12:0] axiRdAddr_15_3_sva;
  reg [7:0] axiRdLen_sva;
  reg [12:0] axiWrAddr_15_3_sva;
  reg select_mask_0_sva;
  reg [63:0] regwr_data_sva;
  reg arb_pick_priority_4_sva;
  reg operator_5_false_operator_5_false_operator_5_false_or_svs;
  reg [2:0] axiRdAddr_2_0_sva_dfm_1;
  reg [2:0] axiWrAddr_2_0_sva_dfm_1;
  reg operator_3_false_2_operator_3_false_2_and_svs_st;
  reg while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st;
  reg while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm;
  reg [7:0] while_else_4_if_if_if_1_for_6_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_47_40_itm_1;
  reg [7:0] while_else_4_if_if_if_1_for_7_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_55_48_itm_1;
  reg [7:0] while_else_4_if_if_if_1_for_8_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_63_56_itm_1;
  reg [63:0] if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0;
  reg [23:0] while_else_4_if_if_axiData_lpi_1_dfm_4_1_63_40;
  reg [7:0] while_else_4_if_if_axiData_lpi_1_dfm_4_1_39_32;
  reg [7:0] while_else_4_if_if_axiData_lpi_1_dfm_4_1_31_24;
  reg [7:0] while_else_4_if_if_axiData_lpi_1_dfm_4_1_23_16;
  reg [7:0] while_else_4_if_if_axiData_lpi_1_dfm_4_1_15_8;
  reg [7:0] while_else_4_if_if_axiData_lpi_1_dfm_4_1_7_0;
  wire if_axi_rd_r_Push_mioi_idat_67_4_mx0c1;
  wire operator_8_false_operator_8_false_nor_mdf_sva_mx1w0;
  wire [63:0] reg_13_sva_dfm_4_mx0w0;
  wire [63:0] reg_12_sva_dfm_4_mx0w0;
  wire [63:0] reg_11_sva_dfm_4_mx0w0;
  wire [63:0] reg_10_sva_dfm_4_mx0w0;
  wire [63:0] reg_9_sva_dfm_4_mx0w0;
  wire [63:0] reg_8_sva_dfm_4_mx0w0;
  wire [63:0] reg_7_sva_dfm_4_mx0w0;
  wire [63:0] reg_6_sva_dfm_4_mx0w0;
  wire [63:0] reg_5_sva_dfm_4_mx0w0;
  wire [63:0] reg_4_sva_dfm_4_mx0w0;
  wire [63:0] reg_3_sva_dfm_4_mx0w0;
  wire [63:0] reg_2_sva_dfm_4_mx0w0;
  wire [63:0] reg_1_sva_dfm_4_mx0w0;
  wire [63:0] reg_0_sva_dfm_4_mx0w0;
  wire [63:0] reg_8_sva_mx1;
  wire [63:0] reg_4_sva_mx1;
  wire [63:0] reg_2_sva_mx1;
  wire [63:0] reg_1_sva_mx1;
  wire [63:0] reg_0_sva_mx1;
  wire [63:0] reg_9_sva_mx1;
  wire [63:0] reg_10_sva_mx1;
  wire [63:0] reg_6_sva_mx1;
  wire [63:0] reg_11_sva_mx1;
  wire [63:0] reg_3_sva_mx1;
  wire [63:0] reg_7_sva_mx1;
  wire [63:0] reg_12_sva_mx1;
  wire [63:0] reg_13_sva_mx1;
  wire [63:0] reg_5_sva_mx1;
  wire operator_5_false_operator_5_false_operator_5_false_or_svs_mx0w0;
  wire while_if_4_while_if_4_and_1_mx0w0;
  wire [2:0] axiRdAddr_2_0_sva_dfm_1_mx1;
  wire [2:0] axiWrAddr_2_0_sva_dfm_1_mx1;
  wire operator_3_false_2_operator_3_false_2_and_svs_st_1_mx0c1;
  wire operator_3_false_3_operator_3_false_3_and_svs_mx0w0;
  wire operator_3_false_2_operator_3_false_2_and_svs_mx0w0;
  wire operator_3_false_1_operator_3_false_1_and_svs_mx0w0;
  wire while_stage_v_2_mx0c1;
  wire while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1_mx0c1;
  wire while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1_mx0c1;
  wire [3:0] operator_17_true_return_1_3_0_sva_mx1;
  wire [12:0] axiRdAddr_15_3_sva_dfm_1_mx0;
  wire [12:0] axiWrAddr_15_3_sva_dfm_1_mx0;
  wire [63:0] axi_rd_resp_data_sva_2;
  wire while_else_4_else_and_13_tmp_1;
  wire while_while_nor_m1c_1;
  wire while_else_4_if_and_14_tmp_1;
  wire while_and_3_m1c_1;
  wire while_else_4_else_and_12_tmp_1;
  wire while_else_4_if_and_13_tmp_1;
  wire while_else_4_else_and_11_tmp_1;
  wire while_else_4_if_and_12_tmp_1;
  wire while_else_4_else_and_10_tmp_1;
  wire while_else_4_if_and_11_tmp_1;
  wire while_else_4_else_and_9_tmp_1;
  wire while_else_4_if_and_10_tmp_1;
  wire while_else_4_else_and_8_tmp_1;
  wire while_else_4_if_and_9_tmp_1;
  wire while_else_4_else_and_7_tmp_1;
  wire while_else_4_else_and_6_tmp_1;
  wire while_else_4_if_and_7_tmp_1;
  wire while_else_4_else_and_5_tmp_1;
  wire while_else_4_if_and_6_tmp_1;
  wire while_else_4_else_and_4_tmp_1;
  wire while_else_4_if_and_5_tmp_1;
  wire while_else_4_else_and_3_tmp_1;
  wire while_else_4_if_and_4_tmp_1;
  wire while_else_4_else_and_2_tmp_1;
  wire while_else_4_if_and_3_tmp_1;
  wire while_else_4_else_and_1_tmp_1;
  wire while_else_4_if_and_2_tmp_1;
  wire while_else_4_else_and_tmp_1;
  wire while_else_4_if_and_1_tmp_1;
  wire [63:0] while_else_4_if_if_if_1_old_data_sva_1;
  wire arb_pick_if_1_not_15;
  wire and_44_rgt;
  wire and_54_rgt;
  wire while_and_rgt;
  wire while_else_4_if_if_regAddr_and_1_cse;
  wire while_else_4_if_if_and_13_cse;
  wire operator_3_false_1_and_cse;
  wire mux_tmp;
  wire mux_tmp_683;
  wire mux_tmp_686;
  wire mux_tmp_687;
  wire nor_tmp_73;
  wire mux_tmp_688;
  wire and_dcpl_141;
  wire nor_tmp_75;
  wire mux_tmp_696;
  wire mux_tmp_697;
  wire mux_tmp_699;
  wire mux_tmp_700;
  wire or_tmp_614;
  wire nand_tmp_110;
  wire mux_tmp_708;
  wire mux_tmp_709;
  wire mux_tmp_712;
  wire mux_tmp_722;
  wire not_tmp_415;
  wire mux_tmp_724;
  wire mux_tmp_730;
  wire not_tmp_422;
  wire mux_tmp_732;
  wire mux_tmp_738;
  wire not_tmp_429;
  wire mux_tmp_740;
  wire mux_tmp_746;
  wire not_tmp_436;
  wire not_tmp_437;
  wire mux_tmp_748;
  wire mux_tmp_754;
  wire not_tmp_445;
  wire mux_tmp_756;
  wire mux_tmp_762;
  wire not_tmp_452;
  wire not_tmp_453;
  wire mux_tmp_764;
  wire mux_tmp_770;
  wire not_tmp_460;
  wire mux_tmp_772;
  wire mux_tmp_778;
  wire not_tmp_468;
  wire mux_tmp_780;
  wire mux_tmp_786;
  wire not_tmp_476;
  wire mux_tmp_788;
  wire or_tmp_728;
  wire mux_tmp_795;
  wire not_tmp_484;
  wire nand_tmp_124;
  wire and_dcpl_196;
  wire nor_tmp_125;
  wire or_tmp_762;
  wire or_tmp_778;
  wire or_tmp_794;
  wire nor_tmp_150;
  wire not_tmp_533;
  wire nor_tmp_158;
  wire nand_198_cse;
  wire nor_151_cse;
  wire or_705_cse;
  wire nand_142_cse_1;
  wire nor_303_cse;
  wire or_735_cse;
  wire and_513_cse;
  wire and_512_cse;
  wire or_927_cse;
  wire and_515_cse;
  wire and_517_cse;
  wire and_499_cse;
  wire and_302_cse;
  wire or_746_cse;
  wire or_841_cse;
  wire or_1037_cse;
  wire mux_833_cse;
  wire mux_884_cse;
  wire and_440_cse;
  wire mux_682_itm;
  wire while_else_4_else_while_else_4_else_and_itm;
  wire while_else_4_if_if_while_else_4_if_if_and_1_itm;
  wire [7:0] while_else_4_if_if_while_else_4_if_if_mux1h_itm;
  wire [7:0] while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm;
  wire [7:0] while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm;
  wire [7:0] while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm;
  wire [7:0] while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm;
  wire [7:0] while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm;
  wire [7:0] while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm;
  wire [7:0] while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm;
  wire mux_683_itm;
  wire mux_684_itm;
  wire mux_725_itm;
  wire mux_730_itm;
  wire mux_738_itm;
  wire mux_746_itm;
  wire mux_754_itm;
  wire mux_762_itm;
  wire mux_770_itm;
  wire mux_778_itm;
  wire mux_786_itm;
  wire mux_794_itm;
  wire [3:0] while_else_4_if_if_regAddr_acc_itm_6_3;
  wire while_if_4_acc_1_itm_16_1;
  wire while_if_4_aelse_acc_itm_16_1;
  wire regwr_addr_and_cse;
  wire while_if_4_and_1_cse;
  wire while_and_110_cse;
  wire while_and_104_cse;
  wire while_and_103_cse;
  wire while_if_4_and_4_cse;

  wire[16:0] while_else_4_if_if_acc_1_nl;
  wire[17:0] nl_while_else_4_if_if_acc_1_nl;
  wire mux_386_nl;
  wire mux_396_nl;
  wire mux_395_nl;
  wire or_344_nl;
  wire mux_394_nl;
  wire or_342_nl;
  wire or_340_nl;
  wire mux_393_nl;
  wire mux_392_nl;
  wire mux_391_nl;
  wire nand_70_nl;
  wire mux_389_nl;
  wire or_337_nl;
  wire mux_384_nl;
  wire mux_383_nl;
  wire nand_68_nl;
  wire nand_67_nl;
  wire mux_382_nl;
  wire mux_403_nl;
  wire mux_402_nl;
  wire mux_401_nl;
  wire or_354_nl;
  wire mux_400_nl;
  wire mux_399_nl;
  wire nand_168_nl;
  wire or_347_nl;
  wire mux_411_nl;
  wire nor_125_nl;
  wire mux_410_nl;
  wire mux_409_nl;
  wire and_354_nl;
  wire mux_406_nl;
  wire and_353_nl;
  wire and_355_nl;
  wire mux_417_nl;
  wire or_376_nl;
  wire mux_416_nl;
  wire nand_75_nl;
  wire mux_415_nl;
  wire mux_414_nl;
  wire mux_687_nl;
  wire mux_686_nl;
  wire and_501_nl;
  wire and_370_nl;
  wire mux_690_nl;
  wire mux_689_nl;
  wire and_503_nl;
  wire and_374_nl;
  wire mux_700_nl;
  wire mux_699_nl;
  wire mux_698_nl;
  wire mux_697_nl;
  wire mux_696_nl;
  wire mux_695_nl;
  wire and_384_nl;
  wire mux_694_nl;
  wire or_710_nl;
  wire and_381_nl;
  wire mux_712_nl;
  wire mux_711_nl;
  wire mux_710_nl;
  wire mux_709_nl;
  wire mux_708_nl;
  wire mux_707_nl;
  wire mux_706_nl;
  wire and_393_nl;
  wire nor_157_nl;
  wire mux_703_nl;
  wire nor_302_nl;
  wire or_720_nl;
  wire mux_726_nl;
  wire and_504_nl;
  wire and_505_nl;
  wire mux_734_nl;
  wire mux_733_nl;
  wire mux_732_nl;
  wire mux_731_nl;
  wire nor_nl;
  wire mux_102_nl;
  wire mux_101_nl;
  wire mux_100_nl;
  wire mux_99_nl;
  wire mux_98_nl;
  wire mux_97_nl;
  wire mux_96_nl;
  wire mux_95_nl;
  wire or_45_nl;
  wire mux_94_nl;
  wire mux_93_nl;
  wire mux_92_nl;
  wire mux_91_nl;
  wire mux_90_nl;
  wire mux_89_nl;
  wire or_74_nl;
  wire mux_742_nl;
  wire mux_741_nl;
  wire mux_740_nl;
  wire mux_739_nl;
  wire nor_387_nl;
  wire mux_126_nl;
  wire mux_125_nl;
  wire mux_124_nl;
  wire mux_123_nl;
  wire mux_122_nl;
  wire mux_121_nl;
  wire mux_120_nl;
  wire or_27_nl;
  wire mux_119_nl;
  wire mux_118_nl;
  wire mux_117_nl;
  wire mux_116_nl;
  wire mux_115_nl;
  wire mux_113_nl;
  wire or_90_nl;
  wire or_121_nl;
  wire mux_750_nl;
  wire mux_749_nl;
  wire mux_748_nl;
  wire mux_747_nl;
  wire and_682_nl;
  wire mux_158_nl;
  wire mux_157_nl;
  wire mux_156_nl;
  wire mux_155_nl;
  wire mux_154_nl;
  wire mux_153_nl;
  wire mux_152_nl;
  wire mux_145_nl;
  wire or_108_nl;
  wire or_120_nl;
  wire mux_150_nl;
  wire mux_142_nl;
  wire mux_141_nl;
  wire mux_140_nl;
  wire mux_139_nl;
  wire and_311_nl;
  wire mux_138_nl;
  wire nor_133_nl;
  wire mux_137_nl;
  wire or_106_nl;
  wire mux_758_nl;
  wire mux_757_nl;
  wire mux_756_nl;
  wire mux_755_nl;
  wire nor_388_nl;
  wire mux_184_nl;
  wire mux_183_nl;
  wire mux_182_nl;
  wire mux_181_nl;
  wire mux_180_nl;
  wire mux_179_nl;
  wire mux_178_nl;
  wire mux_177_nl;
  wire mux_176_nl;
  wire mux_175_nl;
  wire mux_174_nl;
  wire mux_173_nl;
  wire mux_172_nl;
  wire mux_171_nl;
  wire or_134_nl;
  wire mux_766_nl;
  wire mux_765_nl;
  wire mux_764_nl;
  wire mux_763_nl;
  wire nor_389_nl;
  wire mux_210_nl;
  wire mux_209_nl;
  wire mux_208_nl;
  wire mux_207_nl;
  wire mux_206_nl;
  wire mux_205_nl;
  wire mux_204_nl;
  wire mux_203_nl;
  wire mux_202_nl;
  wire mux_201_nl;
  wire mux_200_nl;
  wire mux_199_nl;
  wire mux_198_nl;
  wire mux_197_nl;
  wire or_149_nl;
  wire mux_774_nl;
  wire mux_773_nl;
  wire mux_772_nl;
  wire mux_771_nl;
  wire and_683_nl;
  wire mux_243_nl;
  wire mux_242_nl;
  wire mux_241_nl;
  wire mux_240_nl;
  wire mux_239_nl;
  wire mux_237_nl;
  wire mux_230_nl;
  wire nand_195_nl;
  wire mux_235_nl;
  wire mux_227_nl;
  wire mux_226_nl;
  wire mux_225_nl;
  wire mux_224_nl;
  wire mux_223_nl;
  wire mux_222_nl;
  wire nor_135_nl;
  wire and_318_nl;
  wire or_165_nl;
  wire mux_782_nl;
  wire mux_781_nl;
  wire mux_780_nl;
  wire mux_779_nl;
  wire nor_390_nl;
  wire mux_267_nl;
  wire mux_266_nl;
  wire mux_265_nl;
  wire mux_264_nl;
  wire mux_263_nl;
  wire mux_262_nl;
  wire mux_261_nl;
  wire or_194_nl;
  wire mux_260_nl;
  wire mux_259_nl;
  wire mux_258_nl;
  wire mux_257_nl;
  wire mux_256_nl;
  wire mux_254_nl;
  wire or_192_nl;
  wire mux_790_nl;
  wire mux_789_nl;
  wire mux_788_nl;
  wire mux_787_nl;
  wire nor_391_nl;
  wire mux_293_nl;
  wire mux_292_nl;
  wire mux_291_nl;
  wire mux_290_nl;
  wire mux_289_nl;
  wire mux_288_nl;
  wire mux_287_nl;
  wire mux_286_nl;
  wire mux_285_nl;
  wire mux_284_nl;
  wire mux_283_nl;
  wire mux_282_nl;
  wire mux_281_nl;
  wire mux_280_nl;
  wire nand_143_nl;
  wire mux_798_nl;
  wire mux_797_nl;
  wire mux_796_nl;
  wire mux_795_nl;
  wire nor_392_nl;
  wire mux_319_nl;
  wire mux_318_nl;
  wire mux_317_nl;
  wire mux_316_nl;
  wire mux_315_nl;
  wire mux_314_nl;
  wire mux_313_nl;
  wire mux_312_nl;
  wire mux_311_nl;
  wire mux_310_nl;
  wire mux_309_nl;
  wire mux_308_nl;
  wire mux_307_nl;
  wire mux_306_nl;
  wire or_224_nl;
  wire while_else_4_mux_20_nl;
  wire while_else_4_mux_22_nl;
  wire while_else_4_if_mux_17_nl;
  wire while_if_4_mux1h_3_nl;
  wire while_if_4_while_if_4_or_1_nl;
  wire while_else_4_else_while_else_4_else_or_nl;
  wire while_else_4_if_if_while_else_4_if_if_or_nl;
  wire while_if_4_nand_nl;
  wire mux_808_nl;
  wire mux_807_nl;
  wire nor_305_nl;
  wire mux_806_nl;
  wire and_508_nl;
  wire mux_805_nl;
  wire nor_306_nl;
  wire mux_801_nl;
  wire or_840_nl;
  wire[7:0] while_if_4_else_2_acc_nl;
  wire[8:0] nl_while_if_4_else_2_acc_nl;
  wire mux_505_nl;
  wire mux_504_nl;
  wire nor_129_nl;
  wire and_153_nl;
  wire mux_503_nl;
  wire nor_130_nl;
  wire or_478_nl;
  wire mux_501_nl;
  wire nor_128_nl;
  wire mux_506_nl;
  wire nand_172_nl;
  wire or_486_nl;
  wire mux_550_nl;
  wire mux_549_nl;
  wire and_167_nl;
  wire mux_548_nl;
  wire mux_547_nl;
  wire mux_546_nl;
  wire while_or_25_nl;
  wire while_or_26_nl;
  wire while_and_108_nl;
  wire mux_330_nl;
  wire mux_329_nl;
  wire mux_328_nl;
  wire mux_327_nl;
  wire mux_326_nl;
  wire nor_94_nl;
  wire or_240_nl;
  wire mux_335_nl;
  wire mux_334_nl;
  wire mux_333_nl;
  wire mux_332_nl;
  wire and_323_nl;
  wire mux_331_nl;
  wire nand_144_nl;
  wire and_322_nl;
  wire or_248_nl;
  wire mux_341_nl;
  wire mux_340_nl;
  wire mux_339_nl;
  wire mux_338_nl;
  wire mux_337_nl;
  wire and_307_nl;
  wire mux_336_nl;
  wire nand_140_nl;
  wire or_254_nl;
  wire mux_834_nl;
  wire nand_208_nl;
  wire nand_209_nl;
  wire mux_850_nl;
  wire nand_212_nl;
  wire nand_213_nl;
  wire mux_866_nl;
  wire nand_216_nl;
  wire nand_217_nl;
  wire mux_883_nl;
  wire mux_882_nl;
  wire mux_881_nl;
  wire mux_880_nl;
  wire mux_879_nl;
  wire nor_309_nl;
  wire and_514_nl;
  wire or_940_nl;
  wire and_516_nl;
  wire mux_878_nl;
  wire mux_877_nl;
  wire mux_876_nl;
  wire mux_875_nl;
  wire and_518_nl;
  wire mux_874_nl;
  wire mux_873_nl;
  wire nor_310_nl;
  wire and_520_nl;
  wire mux_872_nl;
  wire mux_871_nl;
  wire mux_870_nl;
  wire and_521_nl;
  wire mux_869_nl;
  wire or_935_nl;
  wire mux_868_nl;
  wire mux_867_nl;
  wire or_1038_nl;
  wire nand_218_nl;
  wire or_930_nl;
  wire and_189_nl;
  wire and_191_nl;
  wire and_193_nl;
  wire and_195_nl;
  wire and_197_nl;
  wire mux_363_nl;
  wire mux_362_nl;
  wire mux_361_nl;
  wire mux_360_nl;
  wire operator_3_false_1_nor_1_nl;
  wire mux_675_nl;
  wire mux_674_nl;
  wire mux_673_nl;
  wire nand_109_nl;
  wire or_602_nl;
  wire mux_672_nl;
  wire mux_671_nl;
  wire or_600_nl;
  wire mux_670_nl;
  wire mux_669_nl;
  wire mux_668_nl;
  wire mux_667_nl;
  wire mux_666_nl;
  wire mux_665_nl;
  wire nand_108_nl;
  wire mux_664_nl;
  wire mux_663_nl;
  wire mux_662_nl;
  wire mux_660_nl;
  wire mux_659_nl;
  wire mux_658_nl;
  wire mux_657_nl;
  wire mux_655_nl;
  wire mux_643_nl;
  wire mux_676_nl;
  wire while_or_13_nl;
  wire while_and_88_nl;
  wire while_and_90_nl;
  wire while_or_12_nl;
  wire while_and_84_nl;
  wire while_and_86_nl;
  wire while_or_11_nl;
  wire while_and_80_nl;
  wire while_and_82_nl;
  wire while_or_10_nl;
  wire while_and_76_nl;
  wire while_and_78_nl;
  wire while_or_9_nl;
  wire while_and_72_nl;
  wire while_and_74_nl;
  wire while_or_8_nl;
  wire while_and_68_nl;
  wire while_and_70_nl;
  wire while_or_7_nl;
  wire while_and_64_nl;
  wire while_and_66_nl;
  wire while_or_6_nl;
  wire while_and_60_nl;
  wire while_and_62_nl;
  wire while_or_5_nl;
  wire while_and_56_nl;
  wire while_and_58_nl;
  wire while_or_4_nl;
  wire while_and_52_nl;
  wire while_and_54_nl;
  wire while_or_3_nl;
  wire while_and_48_nl;
  wire while_and_50_nl;
  wire while_or_2_nl;
  wire while_and_44_nl;
  wire while_and_46_nl;
  wire while_or_1_nl;
  wire while_and_40_nl;
  wire while_and_42_nl;
  wire while_or_15_nl;
  wire while_and_38_nl;
  wire while_and_93_nl;
  wire nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_mux_nl;
  wire while_or_27_nl;
  wire while_or_28_nl;
  wire[6:0] while_else_4_if_if_regAddr_acc_nl;
  wire[8:0] nl_while_else_4_if_if_regAddr_acc_nl;
  wire or_608_nl;
  wire arb_pick_if_1_mux_1_nl;
  wire nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_mux_1_nl;
  wire nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_mux_3_nl;
  wire arb_pick_if_1_mux_3_nl;
  wire[6:0] while_if_4_regAddr_acc_nl;
  wire[8:0] nl_while_if_4_regAddr_acc_nl;
  wire[16:0] while_if_4_acc_1_nl;
  wire[17:0] nl_while_if_4_acc_1_nl;
  wire while_else_4_if_if_and_nl;
  wire while_else_4_if_if_and_1_nl;
  wire while_else_4_if_if_and_4_nl;
  wire while_else_4_if_if_and_5_nl;
  wire while_else_4_if_if_and_6_nl;
  wire while_else_4_if_if_and_7_nl;
  wire while_and_31_nl;
  wire mux_83_nl;
  wire mux_88_nl;
  wire or_661_nl;
  wire mux_109_nl;
  wire mux_114_nl;
  wire nor_137_nl;
  wire mux_133_nl;
  wire or_113_nl;
  wire nand_128_nl;
  wire and_14_nl;
  wire and_13_nl;
  wire mux_148_nl;
  wire mux_165_nl;
  wire mux_170_nl;
  wire nor_139_nl;
  wire mux_191_nl;
  wire mux_196_nl;
  wire or_672_nl;
  wire mux_217_nl;
  wire mux_233_nl;
  wire mux_250_nl;
  wire mux_255_nl;
  wire nor_141_nl;
  wire mux_274_nl;
  wire mux_279_nl;
  wire nor_143_nl;
  wire mux_300_nl;
  wire mux_305_nl;
  wire nor_144_nl;
  wire nor_145_nl;
  wire mux_325_nl;
  wire or_235_nl;
  wire or_293_nl;
  wire nor_106_nl;
  wire mux_371_nl;
  wire and_73_nl;
  wire or_330_nl;
  wire or_690_nl;
  wire or_322_nl;
  wire mux_376_nl;
  wire or_332_nl;
  wire mux_375_nl;
  wire nand_65_nl;
  wire mux_372_nl;
  wire mux_398_nl;
  wire or_351_nl;
  wire and_68_nl;
  wire mux_413_nl;
  wire and_333_nl;
  wire nor_107_nl;
  wire nand_78_nl;
  wire and_107_nl;
  wire mux_426_nl;
  wire mux_425_nl;
  wire and_335_nl;
  wire mux_430_nl;
  wire mux_429_nl;
  wire mux_428_nl;
  wire or_394_nl;
  wire or_391_nl;
  wire mux_435_nl;
  wire mux_434_nl;
  wire nor_110_nl;
  wire mux_454_nl;
  wire mux_453_nl;
  wire mux_957_nl;
  wire nand_88_nl;
  wire mux_450_nl;
  wire mux_685_nl;
  wire mux_447_nl;
  wire mux_445_nl;
  wire mux_444_nl;
  wire mux_443_nl;
  wire and_337_nl;
  wire mux_440_nl;
  wire mux_439_nl;
  wire nand_83_nl;
  wire nand_82_nl;
  wire mux_438_nl;
  wire mux_460_nl;
  wire or_421_nl;
  wire mux_462_nl;
  wire mux_461_nl;
  wire or_418_nl;
  wire or_417_nl;
  wire mux_465_nl;
  wire mux_464_nl;
  wire or_427_nl;
  wire or_426_nl;
  wire or_436_nl;
  wire mux_480_nl;
  wire mux_479_nl;
  wire mux_478_nl;
  wire mux_477_nl;
  wire mux_476_nl;
  wire or_435_nl;
  wire mux_475_nl;
  wire or_434_nl;
  wire mux_468_nl;
  wire mux_467_nl;
  wire mux_466_nl;
  wire and_130_nl;
  wire mux_487_nl;
  wire mux_486_nl;
  wire mux_485_nl;
  wire and_129_nl;
  wire mux_484_nl;
  wire and_127_nl;
  wire mux_483_nl;
  wire and_341_nl;
  wire nor_111_nl;
  wire mux_497_nl;
  wire and_343_nl;
  wire mux_496_nl;
  wire nor_114_nl;
  wire mux_518_nl;
  wire mux_517_nl;
  wire mux_526_nl;
  wire mux_525_nl;
  wire mux_524_nl;
  wire and_161_nl;
  wire mux_528_nl;
  wire mux_523_nl;
  wire mux_522_nl;
  wire mux_521_nl;
  wire mux_520_nl;
  wire mux_537_nl;
  wire mux_544_nl;
  wire mux_543_nl;
  wire and_166_nl;
  wire mux_540_nl;
  wire mux_535_nl;
  wire mux_533_nl;
  wire mux_532_nl;
  wire and_165_nl;
  wire and_164_nl;
  wire mux_531_nl;
  wire and_170_nl;
  wire or_520_nl;
  wire mux_558_nl;
  wire and_171_nl;
  wire or_513_nl;
  wire mux_560_nl;
  wire mux_557_nl;
  wire or_519_nl;
  wire mux_556_nl;
  wire or_515_nl;
  wire mux_567_nl;
  wire mux_574_nl;
  wire mux_573_nl;
  wire nand_97_nl;
  wire mux_570_nl;
  wire mux_565_nl;
  wire mux_563_nl;
  wire or_522_nl;
  wire or_692_nl;
  wire nor_119_nl;
  wire or_581_nl;
  wire mux_613_nl;
  wire mux_612_nl;
  wire and_347_nl;
  wire or_693_nl;
  wire mux_631_nl;
  wire nand_105_nl;
  wire mux_630_nl;
  wire or_593_nl;
  wire mux_629_nl;
  wire or_592_nl;
  wire mux_628_nl;
  wire nor_120_nl;
  wire mux_627_nl;
  wire mux_626_nl;
  wire mux_625_nl;
  wire mux_624_nl;
  wire mux_623_nl;
  wire or_590_nl;
  wire or_588_nl;
  wire mux_621_nl;
  wire mux_620_nl;
  wire mux_619_nl;
  wire mux_618_nl;
  wire mux_617_nl;
  wire mux_616_nl;
  wire mux_615_nl;
  wire nand_164_nl;
  wire mux_640_nl;
  wire mux_639_nl;
  wire mux_638_nl;
  wire mux_651_nl;
  wire mux_680_nl;
  wire mux_679_nl;
  wire mux_677_nl;
  wire nand_89_nl;
  wire mux_457_nl;
  wire mux_456_nl;
  wire nor_123_nl;
  wire mux_578_nl;
  wire mux_577_nl;
  wire or_527_nl;
  wire mux_576_nl;
  wire or_525_nl;
  wire or_524_nl;
  wire mux_582_nl;
  wire mux_581_nl;
  wire mux_580_nl;
  wire mux_579_nl;
  wire nor_131_nl;
  wire mux_589_nl;
  wire mux_588_nl;
  wire or_539_nl;
  wire[16:0] while_if_4_aelse_acc_nl;
  wire[17:0] nl_while_if_4_aelse_acc_nl;
  wire nor_334_nl;
  wire and_572_nl;
  wire nor_335_nl;
  wire and_573_nl;
  wire nor_336_nl;
  wire and_574_nl;
  wire and_380_nl;
  wire and_379_nl;
  wire and_383_nl;
  wire and_382_nl;
  wire nor_338_nl;
  wire and_390_nl;
  wire and_389_nl;
  wire nor_339_nl;
  wire or_722_nl;
  wire and_392_nl;
  wire and_391_nl;
  wire or_730_nl;
  wire or_732_nl;
  wire mux_724_nl;
  wire mux_723_nl;
  wire mux_722_nl;
  wire mux_721_nl;
  wire mux_720_nl;
  wire mux_719_nl;
  wire mux_718_nl;
  wire or_1052_nl;
  wire mux_716_nl;
  wire mux_715_nl;
  wire nand_180_nl;
  wire nor_160_nl;
  wire and_589_nl;
  wire and_590_nl;
  wire nor_343_nl;
  wire nor_344_nl;
  wire and_592_nl;
  wire and_594_nl;
  wire and_595_nl;
  wire nor_345_nl;
  wire nor_346_nl;
  wire and_597_nl;
  wire and_599_nl;
  wire and_600_nl;
  wire nor_347_nl;
  wire nor_348_nl;
  wire and_602_nl;
  wire and_604_nl;
  wire and_605_nl;
  wire nor_349_nl;
  wire nor_350_nl;
  wire and_608_nl;
  wire and_610_nl;
  wire and_611_nl;
  wire nor_351_nl;
  wire nor_352_nl;
  wire and_614_nl;
  wire and_616_nl;
  wire and_617_nl;
  wire nor_353_nl;
  wire nor_354_nl;
  wire and_620_nl;
  wire and_622_nl;
  wire and_623_nl;
  wire nor_355_nl;
  wire nor_356_nl;
  wire and_625_nl;
  wire and_627_nl;
  wire and_628_nl;
  wire and_630_nl;
  wire and_631_nl;
  wire and_632_nl;
  wire and_634_nl;
  wire and_635_nl;
  wire nor_357_nl;
  wire nor_358_nl;
  wire and_637_nl;
  wire mux_799_nl;
  wire and_638_nl;
  wire and_436_nl;
  wire mux_804_nl;
  wire mux_803_nl;
  wire mux_802_nl;
  wire or_849_nl;
  wire mux_832_nl;
  wire mux_831_nl;
  wire mux_830_nl;
  wire mux_829_nl;
  wire mux_828_nl;
  wire nor_367_nl;
  wire or_880_nl;
  wire and_646_nl;
  wire mux_827_nl;
  wire or_879_nl;
  wire mux_826_nl;
  wire mux_825_nl;
  wire and_648_nl;
  wire or_878_nl;
  wire mux_824_nl;
  wire nor_368_nl;
  wire mux_823_nl;
  wire mux_822_nl;
  wire mux_821_nl;
  wire nand_277_nl;
  wire nor_370_nl;
  wire mux_820_nl;
  wire or_1060_nl;
  wire nor_371_nl;
  wire mux_819_nl;
  wire or_872_nl;
  wire or_871_nl;
  wire[17:0] acc_nl;
  wire[18:0] nl_acc_nl;
  wire[15:0] while_else_4_if_if_aelse_mux_2_nl;
  wire while_else_4_if_if_aelse_or_1_nl;
  wire[12:0] while_else_4_if_if_aelse_mux_3_nl;
  wire[2:0] while_else_4_if_if_aelse_while_else_4_if_if_aelse_while_else_4_if_if_aelse_nand_1_nl;
  wire while_else_4_if_if_aelse_not_1_nl;
  wire[12:0] operator_16_false_mux_1_nl;
  wire and_684_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_inst_if_axi_rd_ar_PopNB_mioi_oswt_unreg;
  assign nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_inst_if_axi_rd_ar_PopNB_mioi_oswt_unreg
      = or_dcpl_25 & or_dcpl_3 & or_dcpl_2 & or_234_cse & if_axi_rd_ar_PopNB_mioi_bawt
      & (~ while_asn_25_itm_1) & while_stage_v_1;
  wire  nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_inst_if_axi_wr_aw_PopNB_mioi_oswt_unreg;
  assign nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_inst_if_axi_wr_aw_PopNB_mioi_oswt_unreg
      = and_dcpl_24 & or_dcpl_2 & or_234_cse & if_axi_wr_aw_PopNB_mioi_bawt & (~
      while_asn_30_itm_1) & while_stage_v_1;
  wire  nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_inst_regIn_PopNB_mioi_oswt_unreg;
  assign nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_inst_regIn_PopNB_mioi_oswt_unreg
      = and_dcpl_25 & or_234_cse & regIn_PopNB_mioi_bawt & (~ while_asn_34_itm_1)
      & while_stage_v_1;
  wire  nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_inst_if_axi_rd_r_Push_mioi_oswt_unreg;
  assign nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_inst_if_axi_rd_r_Push_mioi_oswt_unreg
      = while_stage_v_2 & if_axi_rd_r_Push_mioi_bawt & operator_3_false_1_operator_3_false_1_and_svs_st_2;
  wire [70:0] nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_inst_if_axi_rd_r_Push_mioi_idat;
  assign nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_inst_if_axi_rd_r_Push_mioi_idat
      = {if_axi_rd_r_Push_mioi_idat_70 , if_axi_rd_r_Push_mioi_idat_69 , 1'b0 , if_axi_rd_r_Push_mioi_idat_67_4
      , if_axi_rd_r_Push_mioi_idat_3_0};
  wire  nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_inst_if_axi_wr_b_Push_mioi_oswt_unreg;
  assign nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_inst_if_axi_wr_b_Push_mioi_oswt_unreg
      = nor_tmp_25 & while_stage_v_2 & if_axi_wr_b_Push_mioi_bawt & (~ operator_3_false_1_operator_3_false_1_and_svs_st_2);
  wire [5:0] nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_inst_if_axi_wr_b_Push_mioi_idat;
  assign nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_inst_if_axi_wr_b_Push_mioi_idat
      = {if_axi_wr_b_Push_mioi_idat_5 , 1'b0 , if_axi_wr_b_Push_mioi_idat_3_0};
  wire  nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_staller_inst_run_flen_unreg;
  assign nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_staller_inst_run_flen_unreg
      = ~((~((~ while_stage_en_1_mx0w1) & (fsm_output[1]))) | (while_stage_en_1_mx0w1
      & (fsm_output[1])) | (while_stage_v_1 & (~(while_stage_v_2 & or_dcpl_43)) &
      while_or_16_cse_1 & while_or_17_cse_1 & while_or_18_cse_1 & while_or_19_cse_1
      & while_or_cse_1 & while_or_14_cse_1 & (fsm_output[1])) | (while_stage_v_2
      & while_or_cse_1 & while_or_14_cse_1 & (fsm_output[1])));
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_rd_ar_val(if_axi_rd_ar_val),
      .if_axi_rd_ar_rdy(if_axi_rd_ar_rdy),
      .if_axi_rd_ar_msg(if_axi_rd_ar_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_rd_ar_PopNB_mioi_oswt_unreg(nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_ar_PopNB_mioi_inst_if_axi_rd_ar_PopNB_mioi_oswt_unreg),
      .if_axi_rd_ar_PopNB_mioi_bawt(if_axi_rd_ar_PopNB_mioi_bawt),
      .if_axi_rd_ar_PopNB_mioi_iswt0(if_axi_rd_ar_PopNB_mioi_iswt0),
      .if_axi_rd_ar_PopNB_mioi_ivld_mxwt(if_axi_rd_ar_PopNB_mioi_ivld_mxwt),
      .if_axi_rd_ar_PopNB_mioi_idat_mxwt(if_axi_rd_ar_PopNB_mioi_idat_mxwt)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_wr_aw_val(if_axi_wr_aw_val),
      .if_axi_wr_aw_rdy(if_axi_wr_aw_rdy),
      .if_axi_wr_aw_msg(if_axi_wr_aw_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_wr_aw_PopNB_mioi_oswt_unreg(nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_aw_PopNB_mioi_inst_if_axi_wr_aw_PopNB_mioi_oswt_unreg),
      .if_axi_wr_aw_PopNB_mioi_bawt(if_axi_wr_aw_PopNB_mioi_bawt),
      .if_axi_wr_aw_PopNB_mioi_iswt0(if_axi_wr_aw_PopNB_mioi_iswt0),
      .if_axi_wr_aw_PopNB_mioi_ivld_mxwt(if_axi_wr_aw_PopNB_mioi_ivld_mxwt),
      .if_axi_wr_aw_PopNB_mioi_idat_mxwt(if_axi_wr_aw_PopNB_mioi_idat_mxwt)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .regIn_val(regIn_val),
      .regIn_rdy(regIn_rdy),
      .regIn_msg(regIn_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .regIn_PopNB_mioi_oswt_unreg(nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_regIn_PopNB_mioi_inst_regIn_PopNB_mioi_oswt_unreg),
      .regIn_PopNB_mioi_bawt(regIn_PopNB_mioi_bawt),
      .regIn_PopNB_mioi_iswt0(regIn_PopNB_mioi_iswt0),
      .regIn_PopNB_mioi_ivld_mxwt(regIn_PopNB_mioi_ivld_mxwt),
      .regIn_PopNB_mioi_idat_mxwt(regIn_PopNB_mioi_idat_mxwt)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_rd_r_val(if_axi_rd_r_val),
      .if_axi_rd_r_rdy(if_axi_rd_r_rdy),
      .if_axi_rd_r_msg(if_axi_rd_r_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_rd_r_Push_mioi_oswt_unreg(nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_inst_if_axi_rd_r_Push_mioi_oswt_unreg),
      .if_axi_rd_r_Push_mioi_bawt(if_axi_rd_r_Push_mioi_bawt),
      .if_axi_rd_r_Push_mioi_iswt0(if_axi_rd_r_Push_mioi_iswt0),
      .if_axi_rd_r_Push_mioi_wen_comp(if_axi_rd_r_Push_mioi_wen_comp),
      .if_axi_rd_r_Push_mioi_idat(nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_rd_r_Push_mioi_inst_if_axi_rd_r_Push_mioi_idat[70:0])
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_w_PopNB_mioi_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_wr_w_val(if_axi_wr_w_val),
      .if_axi_wr_w_rdy(if_axi_wr_w_rdy),
      .if_axi_wr_w_msg(if_axi_wr_w_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_wr_w_PopNB_mioi_oswt_unreg(and_dcpl_58),
      .if_axi_wr_w_PopNB_mioi_bawt(if_axi_wr_w_PopNB_mioi_bawt),
      .if_axi_wr_w_PopNB_mioi_iswt0(if_axi_wr_w_PopNB_mioi_iswt0),
      .if_axi_wr_w_PopNB_mioi_ivld_mxwt(if_axi_wr_w_PopNB_mioi_ivld_mxwt),
      .if_axi_wr_w_PopNB_mioi_idat_mxwt(if_axi_wr_w_PopNB_mioi_idat_mxwt)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_wr_b_val(if_axi_wr_b_val),
      .if_axi_wr_b_rdy(if_axi_wr_b_rdy),
      .if_axi_wr_b_msg(if_axi_wr_b_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_wr_b_Push_mioi_oswt_unreg(nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_inst_if_axi_wr_b_Push_mioi_oswt_unreg),
      .if_axi_wr_b_Push_mioi_bawt(if_axi_wr_b_Push_mioi_bawt),
      .if_axi_wr_b_Push_mioi_iswt0(if_axi_wr_b_Push_mioi_iswt0),
      .if_axi_wr_b_Push_mioi_wen_comp(if_axi_wr_b_Push_mioi_wen_comp),
      .if_axi_wr_b_Push_mioi_idat(nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_if_axi_wr_b_Push_mioi_inst_if_axi_wr_b_Push_mioi_idat[5:0])
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_staller AxiSlaveToReg2_axi_cfg_standard_14_16_run_staller_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .if_axi_rd_r_Push_mioi_wen_comp(if_axi_rd_r_Push_mioi_wen_comp),
      .if_axi_wr_b_Push_mioi_wen_comp(if_axi_wr_b_Push_mioi_wen_comp),
      .run_flen_unreg(nl_AxiSlaveToReg2_axi_cfg_standard_14_16_run_staller_inst_run_flen_unreg)
    );
  AxiSlaveToReg2_axi_cfg_standard_14_16_run_run_fsm AxiSlaveToReg2_axi_cfg_standard_14_16_run_run_fsm_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign if_axi_wr_bwrite_and_cse = run_wen & (~ (fsm_output[0]));
  assign and_44_rgt = and_dcpl_26 & (~ write_arb_req_sva) & if_axi_wr_w_PopNB_mioi_ivld_mxwt
      & and_dcpl_20 & and_dcpl_19;
  assign and_54_rgt = and_dcpl_26 & (~ read_arb_req_sva) & operator_3_false_1_operator_3_false_1_and_svs_st_1
      & while_stage_v_1;
  assign nor_124_cse = ~(while_if_4_acc_1_itm_16_1 | while_if_4_aelse_acc_itm_16_1);
  assign and_352_cse = (if_axi_wr_w_PopNB_mioi_idat_mxwt[64]) & if_axi_wr_w_PopNB_mioi_ivld_mxwt;
  assign or_310_cse = (while_mux_17_tmp!=8'b00000000);
  assign mux_386_nl = MUX_s_1_2_2(nand_tmp_66, (~ and_tmp_19), arb_next_1_1_sva);
  assign mux_682_itm = MUX_s_1_2_2(mux_tmp_378, mux_386_nl, operator_3_false_3_operator_3_false_3_and_svs_1);
  assign regOut_13_and_cse = run_wen & (~ or_dcpl_43);
  assign nand_198_cse = ~(while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
      & operator_3_false_2_operator_3_false_2_and_svs_st_2);
  assign regOut_8 = reg_regOut_8_cse;
  assign regOut_4 = reg_regOut_4_cse;
  assign or_28_cse = (~ operator_3_false_2_operator_3_false_2_and_svs_st_1) | if_axi_wr_w_PopNB_mioi_bawt;
  assign or_26_cse = (~ operator_3_false_3_operator_3_false_3_and_svs_1) | (while_mux_32_tmp[3]);
  assign nor_151_cse = ~(operator_3_false_2_operator_3_false_2_and_svs_st_1 | (~
      operator_3_false_3_operator_3_false_3_and_svs_1) | (~ operator_3_false_3_operator_3_false_3_and_svs_st_1));
  assign or_705_cse = (~ or_dcpl_2) | (~ while_stage_v_1) | operator_3_false_1_operator_3_false_1_and_svs_1
      | operator_3_false_1_operator_3_false_1_and_svs_st_1;
  assign nor_303_cse = ~(operator_3_false_1_operator_3_false_1_and_svs_2 | (fsm_output[0]));
  assign nand_142_cse_1 = ~(operator_3_false_2_operator_3_false_2_and_svs_st_2 &
      while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
      & while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1 & (~ if_axi_wr_b_Push_mioi_bawt));
  assign and_309_cse = operator_3_false_3_operator_3_false_3_and_svs_1 & (while_mux_32_tmp[3]);
  assign or_735_cse = (~ while_stage_v_1) | operator_3_false_1_operator_3_false_1_and_svs_1;
  assign nor_97_cse = ~((regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (~ (regwr_addr_6_3_sva[2])) | operator_3_false_1_operator_3_false_1_and_svs_2);
  assign or_121_nl = (regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (~ (regwr_addr_6_3_sva[2])) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign mux_151_cse = MUX_s_1_2_2(mux_tmp_144, mux_tmp_143, or_121_nl);
  assign nor_132_cse = ~(nor_97_cse | mux_5_cse);
  assign and_312_cse = (while_mux_32_tmp[1:0]==2'b11);
  assign and_314_cse = (while_else_4_if_if_regAddr_acc_itm_6_3[1:0]==2'b11);
  assign and_499_cse = while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_7_1;
  assign or_210_cse = (while_mux_32_tmp[2:1]!=2'b10);
  assign nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_and_1_cse
      = run_wen & (~(and_256_cse | (fsm_output[0])));
  assign regIn_arb_req_and_cse = run_wen & (and_dcpl_79 | and_dcpl_81);
  assign arb_next_and_cse = run_wen & (~(operator_3_false_operator_3_false_nor_svs_1
      | (~ mux_488_itm) | (fsm_output[0])));
  assign select_mask_and_cse = run_wen & mux_488_itm;
  assign arb_needs_update_and_cse = run_wen & (~((~ mux_489_itm) | (fsm_output[0])));
  assign while_if_4_and_1_cse = (~ operator_3_false_2_operator_3_false_2_and_svs_1)
      & and_dcpl_80;
  assign while_if_4_and_4_cse = if_axi_wr_w_PopNB_mioi_ivld_mxwt & while_and_110_cse;
  assign nor_305_nl = ~(((~(operator_3_false_1_operator_3_false_1_and_svs_st_2 &
      if_axi_rd_r_Push_mioi_bawt)) & while_stage_v_2) | nand_tmp_124);
  assign and_508_nl = operator_3_false_1_operator_3_false_1_and_svs_st_2 & if_axi_rd_r_Push_mioi_bawt;
  assign mux_806_nl = MUX_s_1_2_2(not_tmp_484, mux_tmp_795, and_508_nl);
  assign mux_807_nl = MUX_s_1_2_2(nor_305_nl, mux_806_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign nor_306_nl = ~((~((~ operator_3_false_1_operator_3_false_1_and_svs_st_2)
      | if_axi_rd_r_Push_mioi_bawt | (~ while_stage_v_2))) | nand_tmp_124);
  assign or_840_nl = (~ operator_3_false_1_operator_3_false_1_and_svs_st_2) | if_axi_rd_r_Push_mioi_bawt;
  assign mux_801_nl = MUX_s_1_2_2(not_tmp_484, mux_tmp_795, or_840_nl);
  assign mux_805_nl = MUX_s_1_2_2(nor_306_nl, mux_801_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_808_nl = MUX_s_1_2_2(mux_807_nl, mux_805_nl, nand_142_cse_1);
  assign and_440_cse = mux_808_nl & or_dcpl_2 & or_dcpl_3 & while_stage_v_1 & run_wen;
  assign nor_129_nl = ~(operator_3_false_2_operator_3_false_2_and_svs_1 | (~ nand_tmp_71));
  assign mux_504_nl = MUX_s_1_2_2(nor_129_nl, nand_tmp_71, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign nor_130_nl = ~(if_axi_wr_w_PopNB_mioi_ivld_mxwt | (~ nand_tmp_71));
  assign or_478_nl = operator_3_false_1_operator_3_false_1_and_svs_1 | (~ operator_3_false_2_operator_3_false_2_and_svs_1)
      | (if_axi_wr_w_PopNB_mioi_idat_mxwt[64]);
  assign mux_503_nl = MUX_s_1_2_2(nor_130_nl, nand_tmp_71, or_478_nl);
  assign and_153_nl = if_axi_wr_w_PopNB_mioi_bawt & mux_503_nl;
  assign mux_505_nl = MUX_s_1_2_2(mux_504_nl, and_153_nl, nor_tmp_28);
  assign while_and_rgt = (~ or_dcpl_52) & mux_505_nl & or_dcpl_4 & or_dcpl_3 & or_dcpl_2
      & while_stage_v_1;
  assign operator_3_false_3_and_cse = run_wen & mux_489_itm;
  assign while_and_98_cse = run_wen & (and_dcpl_79 | and_dcpl_81 | or_tmp_576);
  assign while_and_104_cse = operator_3_false_2_operator_3_false_2_and_svs_1 & and_dcpl_81;
  assign while_and_103_cse = (~ operator_3_false_2_operator_3_false_2_and_svs_1)
      & and_dcpl_81;
  assign nor_94_nl = ~(if_axi_rd_r_Push_mioi_bawt | while_nand_2_cse);
  assign mux_326_nl = MUX_s_1_2_2(or_tmp_221, nor_94_nl, or_dcpl_3);
  assign mux_327_nl = MUX_s_1_2_2(or_tmp_221, mux_326_nl, or_dcpl_2);
  assign mux_328_nl = MUX_s_1_2_2(or_tmp_221, mux_327_nl, or_dcpl_4);
  assign mux_329_nl = MUX_s_1_2_2(or_tmp_221, mux_328_nl, and_305_cse);
  assign or_240_nl = (~ while_stage_v_1) | operator_3_false_1_operator_3_false_1_and_svs_st_1;
  assign mux_330_nl = MUX_s_1_2_2(mux_329_nl, or_tmp_221, or_240_nl);
  assign while_else_4_if_if_regAddr_and_1_cse = run_wen & (~ mux_330_nl) & (~ and_dcpl_117);
  assign nand_140_nl = ~((operator_3_false_1_operator_3_false_1_and_svs_2 | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ operator_3_false_2_operator_3_false_2_and_svs_2)) & operator_3_false_2_operator_3_false_2_and_svs_st_2
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
      & while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1 & (~ if_axi_wr_b_Push_mioi_bawt));
  assign mux_336_nl = MUX_s_1_2_2(nand_140_nl, if_axi_rd_r_Push_mioi_bawt, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign and_307_nl = while_stage_v_2 & (~ mux_336_nl);
  assign mux_337_nl = MUX_s_1_2_2(or_tmp_234, and_307_nl, or_dcpl_3);
  assign mux_338_nl = MUX_s_1_2_2(or_tmp_234, mux_337_nl, or_dcpl_2);
  assign mux_339_nl = MUX_s_1_2_2(or_tmp_234, mux_338_nl, or_dcpl_4);
  assign mux_340_nl = MUX_s_1_2_2(or_tmp_234, mux_339_nl, and_305_cse);
  assign or_254_nl = (~ while_stage_v_1) | operator_3_false_1_operator_3_false_1_and_svs_1
      | (~ operator_3_false_2_operator_3_false_2_and_svs_1) | operator_3_false_1_operator_3_false_1_and_svs_st_1;
  assign mux_341_nl = MUX_s_1_2_2(mux_340_nl, or_tmp_234, or_254_nl);
  assign while_else_4_if_if_and_13_cse = run_wen & (~ mux_341_nl) & (~ and_dcpl_117);
  assign and_513_cse = (operator_17_true_return_1_3_0_sva_1[0]) & while_else_4_if_if_for_nor_itm_1;
  assign and_512_cse = (operator_17_true_return_1_3_0_sva_1[2]) & while_else_4_if_if_for_nor_3_itm_1;
  assign or_927_cse = (~ while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1)
      | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1)
      | (~ operator_3_false_2_operator_3_false_2_and_svs_st_2) | if_axi_wr_b_Push_mioi_bawt
      | operator_3_false_1_operator_3_false_1_and_svs_st_2;
  assign and_515_cse = (operator_17_true_return_1_3_0_sva_1[3]) & while_else_4_if_if_for_nor_6_itm_1;
  assign and_517_cse = (operator_17_true_return_1_3_0_sva_1[1]) & while_else_4_if_if_for_nor_1_itm_1;
  assign or_1037_cse = while_else_4_if_if_for_equal_tmp_5_1 | (while_else_4_if_if_regAddr_acc_itm_6_3[3]);
  assign nor_309_nl = ~(while_else_4_if_if_for_equal_tmp_7_1 | while_else_4_if_if_for_equal_tmp_6_1
      | while_else_4_if_if_for_equal_tmp_5_1 | and_512_cse | while_else_4_if_if_for_equal_tmp_12_1
      | while_else_4_if_if_for_equal_tmp_3_1 | and_513_cse | while_else_4_if_if_for_equal_tmp_9_1
      | (while_else_4_if_if_regAddr_acc_itm_6_3[3]) | (~ nor_tmp_150));
  assign and_514_nl = (while_else_4_if_if_regAddr_acc_itm_6_3[3]) & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign mux_879_nl = MUX_s_1_2_2(nor_309_nl, and_514_nl, and_515_cse);
  assign or_940_nl = while_else_4_if_if_for_while_else_4_if_if_for_and_13_itm_1 |
      while_else_4_if_if_for_while_else_4_if_if_for_and_14_itm_1 | while_else_4_if_if_for_equal_tmp_13_1
      | while_else_4_if_if_for_equal_tmp_11_1 | while_else_4_if_if_for_equal_tmp_10_1;
  assign mux_880_nl = MUX_s_1_2_2(mux_879_nl, nor_tmp_158, or_940_nl);
  assign and_516_nl = while_else_4_if_if_for_equal_tmp_10_1 & (while_else_4_if_if_regAddr_acc_itm_6_3[3])
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign mux_881_nl = MUX_s_1_2_2(mux_880_nl, and_516_nl, while_else_4_if_if_regAddr_acc_itm_6_3[1]);
  assign mux_877_nl = MUX_s_1_2_2(not_tmp_533, nor_tmp_150, while_else_4_if_if_for_equal_tmp_10_1);
  assign mux_878_nl = MUX_s_1_2_2(nor_tmp_158, mux_877_nl, while_else_4_if_if_regAddr_acc_itm_6_3[1]);
  assign mux_882_nl = MUX_s_1_2_2(mux_881_nl, mux_878_nl, and_517_cse);
  assign and_518_nl = while_else_4_if_if_for_equal_tmp_9_1 & (while_else_4_if_if_regAddr_acc_itm_6_3[3])
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign mux_874_nl = MUX_s_1_2_2(not_tmp_533, nor_tmp_150, while_else_4_if_if_for_equal_tmp_9_1);
  assign mux_875_nl = MUX_s_1_2_2(and_518_nl, mux_874_nl, and_513_cse);
  assign nor_310_nl = ~((~ while_else_4_if_if_for_equal_tmp_3_1) | (while_else_4_if_if_regAddr_acc_itm_6_3[3])
      | (~ nor_tmp_150));
  assign and_520_nl = (while_else_4_if_if_for_equal_tmp_3_1 | (while_else_4_if_if_regAddr_acc_itm_6_3[3]))
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign mux_873_nl = MUX_s_1_2_2(nor_310_nl, and_520_nl, while_else_4_if_if_for_equal_tmp_11_1);
  assign mux_876_nl = MUX_s_1_2_2(mux_875_nl, mux_873_nl, while_else_4_if_if_regAddr_acc_itm_6_3[1]);
  assign mux_883_nl = MUX_s_1_2_2(mux_882_nl, mux_876_nl, while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign and_521_nl = while_else_4_if_if_for_equal_tmp_12_1 & (while_else_4_if_if_regAddr_acc_itm_6_3[3])
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign mux_869_nl = MUX_s_1_2_2(not_tmp_533, nor_tmp_150, while_else_4_if_if_for_equal_tmp_12_1);
  assign mux_870_nl = MUX_s_1_2_2(and_521_nl, mux_869_nl, and_512_cse);
  assign or_935_nl = (~ while_else_4_if_if_for_equal_tmp_6_1) | (while_else_4_if_if_regAddr_acc_itm_6_3[3])
      | (~ nor_tmp_150);
  assign mux_871_nl = MUX_s_1_2_2((~ mux_870_nl), or_935_nl, while_else_4_if_if_regAddr_acc_itm_6_3[1]);
  assign or_1038_nl = (~ while_else_4_if_if_for_equal_tmp_5_1) | (while_else_4_if_if_regAddr_acc_itm_6_3[3])
      | (~ nor_tmp_150);
  assign nand_218_nl = ~(or_1037_cse & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1);
  assign mux_867_nl = MUX_s_1_2_2(or_1038_nl, nand_218_nl, while_else_4_if_if_for_equal_tmp_13_1);
  assign or_930_nl = (~ while_else_4_if_if_for_equal_tmp_7_1) | (while_else_4_if_if_regAddr_acc_itm_6_3[3])
      | (~ nor_tmp_150);
  assign mux_868_nl = MUX_s_1_2_2(mux_867_nl, or_930_nl, while_else_4_if_if_regAddr_acc_itm_6_3[1]);
  assign mux_872_nl = MUX_s_1_2_2(mux_871_nl, mux_868_nl, while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign mux_884_cse = MUX_s_1_2_2((~ mux_883_nl), mux_872_nl, while_else_4_if_if_regAddr_acc_itm_6_3[2]);
  assign operator_3_false_2_and_2_cse = run_wen & (~((~ and_dcpl_26) | and_dcpl_83
      | (~ while_stage_v_1)));
  assign operator_3_false_1_nor_1_nl = ~(or_dcpl_4 | (~ or_dcpl_17));
  assign mux_360_nl = MUX_s_1_2_2(or_dcpl_17, operator_3_false_1_nor_1_nl, or_dcpl_3);
  assign mux_361_nl = MUX_s_1_2_2(or_dcpl_17, mux_360_nl, or_dcpl_2);
  assign mux_362_nl = MUX_s_1_2_2(or_dcpl_17, mux_361_nl, or_234_cse);
  assign mux_363_nl = MUX_s_1_2_2(or_dcpl_17, mux_362_nl, while_stage_v_1);
  assign operator_3_false_1_and_cse = ~((~ run_wen) | mux_363_nl | and_dcpl_35);
  assign regwr_addr_and_cse = run_wen & (~((~ and_dcpl_26) | and_dcpl_83 | regIn_arb_req_sva
      | (~ while_stage_v_1)));
  assign operator_8_false_operator_8_false_nor_mdf_sva_mx1w0 = ~((axiRdLen_sva_dfm_1_mx0!=8'b00000000));
  assign while_or_13_nl = ((~ while_else_4_else_and_13_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_14_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_88_nl = while_else_4_else_and_13_tmp_1 & while_while_nor_m1c_1;
  assign while_and_90_nl = while_else_4_if_and_14_tmp_1 & while_and_3_m1c_1;
  assign reg_13_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_13_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_13_nl
      , while_and_88_nl , while_and_90_nl});
  assign while_or_12_nl = ((~ while_else_4_else_and_12_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_13_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_84_nl = while_else_4_else_and_12_tmp_1 & while_while_nor_m1c_1;
  assign while_and_86_nl = while_else_4_if_and_13_tmp_1 & while_and_3_m1c_1;
  assign reg_12_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_12_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_12_nl
      , while_and_84_nl , while_and_86_nl});
  assign while_or_11_nl = ((~ while_else_4_else_and_11_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_12_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_80_nl = while_else_4_else_and_11_tmp_1 & while_while_nor_m1c_1;
  assign while_and_82_nl = while_else_4_if_and_12_tmp_1 & while_and_3_m1c_1;
  assign reg_11_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_11_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_11_nl
      , while_and_80_nl , while_and_82_nl});
  assign while_or_10_nl = ((~ while_else_4_else_and_10_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_11_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_76_nl = while_else_4_else_and_10_tmp_1 & while_while_nor_m1c_1;
  assign while_and_78_nl = while_else_4_if_and_11_tmp_1 & while_and_3_m1c_1;
  assign reg_10_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_10_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_10_nl
      , while_and_76_nl , while_and_78_nl});
  assign while_or_9_nl = ((~ while_else_4_else_and_9_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_10_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_72_nl = while_else_4_else_and_9_tmp_1 & while_while_nor_m1c_1;
  assign while_and_74_nl = while_else_4_if_and_10_tmp_1 & while_and_3_m1c_1;
  assign reg_9_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_9_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_9_nl
      , while_and_72_nl , while_and_74_nl});
  assign while_or_8_nl = ((~ while_else_4_else_and_8_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_9_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_68_nl = while_else_4_else_and_8_tmp_1 & while_while_nor_m1c_1;
  assign while_and_70_nl = while_else_4_if_and_9_tmp_1 & while_and_3_m1c_1;
  assign reg_8_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_regOut_8_cse, regwr_data_sva,
      ({while_else_4_if_if_while_else_4_if_if_mux1h_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_8_nl
      , while_and_68_nl , while_and_70_nl});
  assign while_or_7_nl = ((~ while_else_4_else_and_7_tmp_1) & while_while_nor_m1c_1)
      | ((~ and_499_cse) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_64_nl = while_else_4_else_and_7_tmp_1 & while_while_nor_m1c_1;
  assign while_and_66_nl = and_499_cse & while_and_3_m1c_1;
  assign reg_7_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_7_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_7_nl
      , while_and_64_nl , while_and_66_nl});
  assign while_or_6_nl = ((~ while_else_4_else_and_6_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_7_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_60_nl = while_else_4_else_and_6_tmp_1 & while_while_nor_m1c_1;
  assign while_and_62_nl = while_else_4_if_and_7_tmp_1 & while_and_3_m1c_1;
  assign reg_6_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_6_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_6_nl
      , while_and_60_nl , while_and_62_nl});
  assign while_or_5_nl = ((~ while_else_4_else_and_5_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_6_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_56_nl = while_else_4_else_and_5_tmp_1 & while_while_nor_m1c_1;
  assign while_and_58_nl = while_else_4_if_and_6_tmp_1 & while_and_3_m1c_1;
  assign reg_5_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_5_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_5_nl
      , while_and_56_nl , while_and_58_nl});
  assign while_or_4_nl = ((~ while_else_4_else_and_4_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_5_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_52_nl = while_else_4_else_and_4_tmp_1 & while_while_nor_m1c_1;
  assign while_and_54_nl = while_else_4_if_and_5_tmp_1 & while_and_3_m1c_1;
  assign reg_4_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_regOut_4_cse, regwr_data_sva,
      ({while_else_4_if_if_while_else_4_if_if_mux1h_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_4_nl
      , while_and_52_nl , while_and_54_nl});
  assign while_or_3_nl = ((~ while_else_4_else_and_3_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_4_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_48_nl = while_else_4_else_and_3_tmp_1 & while_while_nor_m1c_1;
  assign while_and_50_nl = while_else_4_if_and_4_tmp_1 & while_and_3_m1c_1;
  assign reg_3_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_3_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_3_nl
      , while_and_48_nl , while_and_50_nl});
  assign while_or_2_nl = ((~ while_else_4_else_and_2_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_3_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_44_nl = while_else_4_else_and_2_tmp_1 & while_while_nor_m1c_1;
  assign while_and_46_nl = while_else_4_if_and_3_tmp_1 & while_and_3_m1c_1;
  assign reg_2_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_2_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_2_nl
      , while_and_44_nl , while_and_46_nl});
  assign while_or_1_nl = ((~ while_else_4_else_and_1_tmp_1) & while_while_nor_m1c_1)
      | ((~ while_else_4_if_and_2_tmp_1) & while_and_3_m1c_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign while_and_40_nl = while_else_4_else_and_1_tmp_1 & while_while_nor_m1c_1;
  assign while_and_42_nl = while_else_4_if_and_2_tmp_1 & while_and_3_m1c_1;
  assign reg_1_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_1_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_1_nl
      , while_and_40_nl , while_and_42_nl});
  assign while_or_15_nl = ((~ while_else_4_else_and_tmp_1) & while_while_nor_m1c_1)
      | operator_3_false_1_operator_3_false_1_and_svs_2 | ((~ while_else_4_if_and_1_tmp_1)
      & while_and_3_m1c_1);
  assign while_and_38_nl = while_else_4_else_and_tmp_1 & while_while_nor_m1c_1;
  assign while_and_93_nl = while_else_4_if_and_1_tmp_1 & while_and_3_m1c_1;
  assign reg_0_sva_dfm_4_mx0w0 = MUX1HOT_v_64_3_2(reg_0_sva, regwr_data_sva, ({while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm
      , while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm}), {while_or_15_nl
      , while_and_38_nl , while_and_93_nl});
  assign while_stage_en_1_mx0w1 = while_or_16_cse_1 & while_or_17_cse_1 & while_or_18_cse_1
      & while_or_19_cse_1 & while_or_cse_1 & while_or_14_cse_1;
  assign reg_8_sva_mx1 = MUX_v_64_2_2(reg_regOut_8_cse, reg_8_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_4_sva_mx1 = MUX_v_64_2_2(reg_regOut_4_cse, reg_4_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_2_sva_mx1 = MUX_v_64_2_2(reg_2_sva, reg_2_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_1_sva_mx1 = MUX_v_64_2_2(reg_1_sva, reg_1_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_0_sva_mx1 = MUX_v_64_2_2(reg_0_sva, reg_0_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_9_sva_mx1 = MUX_v_64_2_2(reg_9_sva, reg_9_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_10_sva_mx1 = MUX_v_64_2_2(reg_10_sva, reg_10_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_6_sva_mx1 = MUX_v_64_2_2(reg_6_sva, reg_6_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_11_sva_mx1 = MUX_v_64_2_2(reg_11_sva, reg_11_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_3_sva_mx1 = MUX_v_64_2_2(reg_3_sva, reg_3_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_7_sva_mx1 = MUX_v_64_2_2(reg_7_sva, reg_7_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_12_sva_mx1 = MUX_v_64_2_2(reg_12_sva, reg_12_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_13_sva_mx1 = MUX_v_64_2_2(reg_13_sva, reg_13_sva_dfm_4_mx0w0, while_stage_v_2);
  assign reg_5_sva_mx1 = MUX_v_64_2_2(reg_5_sva, reg_5_sva_dfm_4_mx0w0, while_stage_v_2);
  assign nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_mux_nl
      = MUX_s_1_2_2(regIn_arb_req_sva_mx1, arb_pick_priority_3_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1);
  assign nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm_mx0w0
      = nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_mux_nl
      & (~ arb_pick_priority_4_sva_mx0w0);
  assign nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm_mx0w0
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1 & (~ arb_pick_priority_4_sva_mx0w0);
  assign arb_pick_if_1_and_tmp_2_mx0w0 = (~ nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm_mx0w0)
      & nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm_mx0w0;
  assign arb_pick_if_1_and_stg_1_0_mx0w0 = ~(nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm_mx0w0
      | nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm_mx0w0);
  assign arb_pick_priority_4_sva_mx0w0 = arb_next_1_2_sva & regIn_arb_req_sva_mx1;
  assign arb_pick_priority_4_sva_mx1 = MUX_s_1_2_2(arb_pick_priority_4_sva, arb_pick_priority_4_sva_mx0w0,
      mux_481_itm);
  assign operator_5_false_operator_5_false_operator_5_false_or_svs_mx0w0 = read_arb_req_sva_mx1
      | regIn_arb_req_sva_mx1 | write_arb_req_sva_mx1;
  assign operator_5_false_operator_5_false_operator_5_false_or_svs_mx1 = MUX_s_1_2_2(operator_5_false_operator_5_false_operator_5_false_or_svs,
      operator_5_false_operator_5_false_operator_5_false_or_svs_mx0w0, mux_481_itm);
  assign while_else_4_else_while_else_4_else_and_itm = while_while_or_2_tmp & (~
      operator_3_false_3_operator_3_false_3_and_svs_1);
  assign while_and_110_cse = operator_3_false_2_operator_3_false_2_and_svs_1 & and_dcpl_80;
  assign while_or_27_nl = and_dcpl_77 | while_and_110_cse;
  assign regIn_arb_req_sva_mx1 = MUX1HOT_s_1_3_2(while_while_or_2_tmp, while_else_4_else_while_else_4_else_and_itm,
      regIn_arb_req_sva, {while_or_27_nl , while_if_4_and_1_cse , (~ while_stage_v_1)});
  assign while_if_4_while_if_4_and_1_mx0w0 = while_while_or_tmp & (~ operator_8_false_operator_8_false_nor_mdf_sva_mx1);
  assign read_arb_req_sva_mx1 = MUX1HOT_s_1_3_2(while_if_4_while_if_4_and_1_mx0w0,
      while_while_or_tmp, read_arb_req_sva, {and_dcpl_77 , and_dcpl_80 , (~ while_stage_v_1)});
  assign while_else_4_if_if_while_else_4_if_if_and_1_itm = while_while_or_1_tmp &
      (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[64]));
  assign while_or_28_nl = and_dcpl_77 | while_if_4_and_1_cse | ((~ if_axi_wr_w_PopNB_mioi_ivld_mxwt)
      & while_and_110_cse);
  assign write_arb_req_sva_mx1 = MUX1HOT_s_1_3_2(while_while_or_1_tmp, while_else_4_if_if_while_else_4_if_if_and_1_itm,
      write_arb_req_sva, {while_or_28_nl , while_if_4_and_4_cse , (~ while_stage_v_1)});
  assign axiRdAddr_2_0_sva_dfm_1_mx1 = MUX_v_3_2_2((if_axi_rd_ar_PopNB_mioi_idat_mxwt[6:4]),
      axiRdAddr_2_0_sva_dfm_1, or_dcpl_51);
  assign axiWrAddr_2_0_sva_dfm_1_mx1 = MUX_v_3_2_2((if_axi_wr_aw_PopNB_mioi_idat_mxwt[6:4]),
      axiWrAddr_2_0_sva_dfm_1, or_dcpl_52);
  assign operator_8_false_operator_8_false_nor_mdf_sva_mx1 = MUX_s_1_2_2(operator_8_false_operator_8_false_nor_mdf_sva,
      operator_8_false_operator_8_false_nor_mdf_sva_mx1w0, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign operator_3_false_3_operator_3_false_3_and_svs_mx0w0 = select_mask_2_1_sva_dfm_1_mx0
      & (~(select_mask_2_1_sva_dfm_0_mx0 | select_mask_0_sva_dfm_mx0));
  assign operator_3_false_2_operator_3_false_2_and_svs_mx0w0 = select_mask_2_1_sva_dfm_0_mx0
      & (~(select_mask_2_1_sva_dfm_1_mx0 | select_mask_0_sva_dfm_mx0));
  assign operator_3_false_1_operator_3_false_1_and_svs_mx0w0 = select_mask_0_sva_dfm_mx0
      & (~(select_mask_2_1_sva_dfm_1_mx0 | select_mask_2_1_sva_dfm_0_mx0));
  assign nl_while_else_4_if_if_regAddr_acc_nl = ({(axiWrAddr_15_3_sva_dfm_1_mx0[3:0])
      , axiWrAddr_2_0_sva_dfm_1_mx1}) - (baseAddr[6:0]);
  assign while_else_4_if_if_regAddr_acc_nl = nl_while_else_4_if_if_regAddr_acc_nl[6:0];
  assign while_else_4_if_if_regAddr_acc_itm_6_3 = readslicef_7_4_3(while_else_4_if_if_regAddr_acc_nl);
  assign or_608_nl = (~(if_axi_wr_w_PopNB_mioi_ivld_mxwt & operator_3_false_2_operator_3_false_2_and_svs_st_1))
      | operator_3_false_1_operator_3_false_1_and_svs_st_1;
  assign operator_17_true_return_1_3_0_sva_mx1 = MUX_v_4_2_2(while_else_4_if_if_regAddr_acc_itm_6_3,
      operator_17_true_return_1_3_0_sva_1, or_608_nl);
  assign select_mask_2_1_sva_dfm_0_mx0 = MUX_s_1_2_2(arb_pick_return_2_1_lpi_1_dfm_1_0_1,
      select_mask_2_1_sva_0, and_dcpl_130);
  assign select_mask_2_1_sva_dfm_1_mx0 = MUX_s_1_2_2(arb_pick_return_2_1_lpi_1_dfm_1_1_1,
      select_mask_2_1_sva_1, and_dcpl_130);
  assign select_mask_0_sva_dfm_mx0 = MUX_s_1_2_2(arb_pick_return_0_lpi_1_dfm_2, select_mask_0_sva,
      and_dcpl_130);
  assign nvhls_set_slc_Arbiter_3U_Roundrobin_Mask_nvhls_nvhls_t_2U_nvuint_t_X_temp_2_1_sva_1_1
      = arb_pick_priority_4_sva_mx0w0 | (nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm_mx0w0
      & (~ nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm_mx0w0));
  assign arb_pick_priority_3_sva_1 = arb_next_1_1_sva & write_arb_req_sva_mx1;
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1 = arb_pick_priority_3_sva_1
      | read_arb_req_sva_mx1;
  assign arb_pick_if_1_mux_1_nl = MUX_s_1_2_2(arb_pick_if_1_and_tmp_2, arb_pick_if_1_and_tmp_2_mx0w0,
      mux_481_itm);
  assign arb_pick_return_0_lpi_1_dfm_2 = arb_pick_if_1_mux_1_nl & operator_5_false_operator_5_false_operator_5_false_or_svs_mx1
      & (~ operator_3_false_operator_3_false_nor_svs_1);
  assign arb_pick_return_2_1_lpi_1_dfm_1_1_1 = nvhls_set_slc_Arbiter_3U_Roundrobin_Mask_nvhls_nvhls_t_2U_nvuint_t_X_temp_2_1_sva_1_1
      & operator_5_false_operator_5_false_operator_5_false_or_svs_mx1;
  assign nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_mux_1_nl
      = MUX_s_1_2_2(nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm,
      nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm_mx0w0,
      mux_481_itm);
  assign nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_mux_3_nl
      = MUX_s_1_2_2(nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm,
      nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm_mx0w0,
      mux_481_itm);
  assign arb_pick_if_1_mux_3_nl = MUX_s_1_2_2(arb_pick_if_1_and_stg_1_0, arb_pick_if_1_and_stg_1_0_mx0w0,
      mux_481_itm);
  assign arb_pick_return_2_1_lpi_1_dfm_1_0_1 = ((nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_mux_1_nl
      & nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_mux_3_nl
      & (~ arb_pick_priority_4_sva_mx1)) | (arb_pick_if_1_mux_3_nl & (~ arb_pick_priority_4_sva_mx1)))
      & operator_5_false_operator_5_false_operator_5_false_or_svs_mx1 & (~ operator_3_false_operator_3_false_nor_svs_1);
  assign operator_3_false_operator_3_false_nor_svs_1 = ~(regIn_arb_req_sva_mx1 |
      write_arb_req_sva_mx1 | read_arb_req_sva_mx1);
  assign axiRdAddr_15_3_sva_dfm_1_mx0 = MUX_v_13_2_2((if_axi_rd_ar_PopNB_mioi_idat_mxwt[19:7]),
      axiRdAddr_15_3_sva, or_dcpl_51);
  assign axiRdLen_sva_dfm_1_mx0 = MUX_v_8_2_2((if_axi_rd_ar_PopNB_mioi_idat_mxwt[27:20]),
      axiRdLen_sva, or_dcpl_51);
  assign axiWrAddr_15_3_sva_dfm_1_mx0 = MUX_v_13_2_2((if_axi_wr_aw_PopNB_mioi_idat_mxwt[19:7]),
      axiWrAddr_15_3_sva, or_dcpl_52);
  assign nl_while_if_4_regAddr_acc_nl = ({(axiRdAddr_15_3_sva_dfm_1_mx0[3:0]) , axiRdAddr_2_0_sva_dfm_1_mx1})
      - (baseAddr[6:0]);
  assign while_if_4_regAddr_acc_nl = nl_while_if_4_regAddr_acc_nl[6:0];
  assign axi_rd_resp_data_sva_2 = MUX_v_64_14_2(reg_0_sva_mx1, reg_1_sva_mx1, reg_2_sva_mx1,
      reg_3_sva_mx1, reg_4_sva_mx1, reg_5_sva_mx1, reg_6_sva_mx1, reg_7_sva_mx1,
      reg_8_sva_mx1, reg_9_sva_mx1, reg_10_sva_mx1, reg_11_sva_mx1, reg_12_sva_mx1,
      reg_13_sva_mx1, readslicef_7_4_3(while_if_4_regAddr_acc_nl));
  assign nl_while_if_4_acc_1_nl = ({1'b1 , axiRdAddr_15_3_sva_dfm_1_mx0 , axiRdAddr_2_0_sva_dfm_1_mx1})
      + conv_u2u_16_17(~ baseAddr) + 17'b00000000000000001;
  assign while_if_4_acc_1_nl = nl_while_if_4_acc_1_nl[16:0];
  assign while_if_4_acc_1_itm_16_1 = readslicef_17_1_16(while_if_4_acc_1_nl);
  assign while_while_or_1_tmp = if_axi_wr_aw_PopNB_mioi_ivld_mxwt | write_arb_req_sva;
  assign while_while_or_2_tmp = regIn_PopNB_mioi_ivld_mxwt | regIn_arb_req_sva;
  assign while_while_or_tmp = if_axi_rd_ar_PopNB_mioi_ivld_mxwt | read_arb_req_sva;
  assign while_else_4_if_if_and_nl = (~ (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[2]))
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign while_else_4_if_if_and_1_nl = (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[2])
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign while_else_4_if_if_while_else_4_if_if_mux1h_itm = MUX1HOT_v_8_3_2((if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0[63:56]),
      while_else_4_if_if_if_1_for_8_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_63_56_itm_1,
      (while_else_4_if_if_axiData_lpi_1_dfm_4_1_63_40[23:16]), {(~ while_else_4_if_if_while_else_4_if_if_nand_tmp_1)
      , while_else_4_if_if_and_nl , while_else_4_if_if_and_1_nl});
  assign while_else_4_if_if_and_4_nl = (~ (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[1]))
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign while_else_4_if_if_and_5_nl = (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[1])
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_itm
      = MUX1HOT_v_8_3_2((if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0[55:48]), while_else_4_if_if_if_1_for_7_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_55_48_itm_1,
      (while_else_4_if_if_axiData_lpi_1_dfm_4_1_63_40[15:8]), {(~ while_else_4_if_if_while_else_4_if_if_nand_tmp_1)
      , while_else_4_if_if_and_4_nl , while_else_4_if_if_and_5_nl});
  assign while_else_4_if_if_and_6_nl = (~ (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[0]))
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign while_else_4_if_if_and_7_nl = (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[0])
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux1h_1_itm
      = MUX1HOT_v_8_3_2((if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0[47:40]), while_else_4_if_if_if_1_for_6_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_47_40_itm_1,
      (while_else_4_if_if_axiData_lpi_1_dfm_4_1_63_40[7:0]), {(~ while_else_4_if_if_while_else_4_if_if_nand_tmp_1)
      , while_else_4_if_if_and_6_nl , while_else_4_if_if_and_7_nl});
  assign while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_2_itm = MUX_v_8_2_2((if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0[39:32]),
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_39_32, while_else_4_if_if_while_else_4_if_if_nand_tmp_1);
  assign while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_3_itm = MUX_v_8_2_2((if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0[31:24]),
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_31_24, while_else_4_if_if_while_else_4_if_if_nand_tmp_1);
  assign while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_4_itm = MUX_v_8_2_2((if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0[23:16]),
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_23_16, while_else_4_if_if_while_else_4_if_if_nand_tmp_1);
  assign while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_5_itm = MUX_v_8_2_2((if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0[15:8]),
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_15_8, while_else_4_if_if_while_else_4_if_if_nand_tmp_1);
  assign while_else_4_if_if_while_else_4_if_if_while_else_4_if_if_mux_6_itm = MUX_v_8_2_2((if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0[7:0]),
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_7_0, while_else_4_if_if_while_else_4_if_if_nand_tmp_1);
  assign while_else_4_else_if_and_stg_2_0_sva_1 = while_else_4_else_if_and_stg_1_0_sva_1
      & (~ (regwr_addr_6_3_sva[2]));
  assign while_else_4_else_if_and_stg_2_1_sva_1 = while_else_4_else_if_and_stg_1_1_sva_1
      & (~ (regwr_addr_6_3_sva[2]));
  assign while_else_4_else_if_and_stg_2_2_sva_1 = while_else_4_else_if_and_stg_1_2_sva_1
      & (~ (regwr_addr_6_3_sva[2]));
  assign while_else_4_else_if_and_stg_1_2_sva_1 = (regwr_addr_6_3_sva[1:0]==2'b10);
  assign while_else_4_else_if_and_stg_2_3_sva_1 = while_else_4_else_if_and_stg_1_3_sva_1
      & (~ (regwr_addr_6_3_sva[2]));
  assign while_else_4_else_if_and_stg_1_3_sva_1 = (regwr_addr_6_3_sva[1:0]==2'b11);
  assign while_else_4_else_if_and_stg_2_4_sva_1 = while_else_4_else_if_and_stg_1_0_sva_1
      & (regwr_addr_6_3_sva[2]);
  assign while_else_4_else_if_and_stg_2_5_sva_1 = while_else_4_else_if_and_stg_1_1_sva_1
      & (regwr_addr_6_3_sva[2]);
  assign while_else_4_else_if_and_stg_1_0_sva_1 = ~((regwr_addr_6_3_sva[1:0]!=2'b00));
  assign while_else_4_else_if_and_stg_1_1_sva_1 = (regwr_addr_6_3_sva[1:0]==2'b01);
  assign while_else_4_else_and_13_tmp_1 = while_else_4_else_if_and_stg_2_5_sva_1
      & (regwr_addr_6_3_sva[3]) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_while_nor_m1c_1 = ~(operator_3_false_2_operator_3_false_2_and_svs_2
      | operator_3_false_1_operator_3_false_1_and_svs_2);
  assign while_else_4_if_and_14_tmp_1 = while_else_4_if_if_for_equal_tmp_13_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_3_m1c_1 = operator_3_false_2_operator_3_false_2_and_svs_2 & (~
      operator_3_false_1_operator_3_false_1_and_svs_2);
  assign while_else_4_else_and_12_tmp_1 = while_else_4_else_if_and_stg_2_4_sva_1
      & (regwr_addr_6_3_sva[3]) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_13_tmp_1 = while_else_4_if_if_for_equal_tmp_12_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_11_tmp_1 = while_else_4_else_if_and_stg_2_3_sva_1
      & (regwr_addr_6_3_sva[3]) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_12_tmp_1 = while_else_4_if_if_for_equal_tmp_11_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_10_tmp_1 = while_else_4_else_if_and_stg_2_2_sva_1
      & (regwr_addr_6_3_sva[3]) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_11_tmp_1 = while_else_4_if_if_for_equal_tmp_10_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_9_tmp_1 = while_else_4_else_if_and_stg_2_1_sva_1 &
      (regwr_addr_6_3_sva[3]) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_10_tmp_1 = while_else_4_if_if_for_equal_tmp_9_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_8_tmp_1 = while_else_4_else_if_and_stg_2_0_sva_1 &
      (regwr_addr_6_3_sva[3]) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_9_tmp_1 = and_515_cse & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_7_tmp_1 = while_else_4_else_if_and_stg_1_3_sva_1 &
      (regwr_addr_6_3_sva[3:2]==2'b01) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_else_and_6_tmp_1 = while_else_4_else_if_and_stg_1_2_sva_1 &
      (regwr_addr_6_3_sva[3:2]==2'b01) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_7_tmp_1 = while_else_4_if_if_for_equal_tmp_6_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_5_tmp_1 = while_else_4_else_if_and_stg_2_5_sva_1 &
      (~ (regwr_addr_6_3_sva[3])) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_6_tmp_1 = while_else_4_if_if_for_equal_tmp_5_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_4_tmp_1 = while_else_4_else_if_and_stg_2_4_sva_1 &
      (~ (regwr_addr_6_3_sva[3])) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_5_tmp_1 = and_512_cse & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_3_tmp_1 = while_else_4_else_if_and_stg_2_3_sva_1 &
      (~ (regwr_addr_6_3_sva[3])) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_4_tmp_1 = while_else_4_if_if_for_equal_tmp_3_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_2_tmp_1 = while_else_4_else_if_and_stg_2_2_sva_1 &
      (~ (regwr_addr_6_3_sva[3])) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_3_tmp_1 = and_517_cse & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_1_tmp_1 = while_else_4_else_if_and_stg_2_1_sva_1 &
      (~ (regwr_addr_6_3_sva[3])) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_2_tmp_1 = and_513_cse & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_else_4_else_and_tmp_1 = while_else_4_else_if_and_stg_2_0_sva_1 & (~
      (regwr_addr_6_3_sva[3])) & operator_3_false_3_operator_3_false_3_and_svs_2;
  assign while_else_4_if_and_1_tmp_1 = (~(and_513_cse | and_517_cse | while_else_4_if_if_for_equal_tmp_3_1
      | and_512_cse | while_else_4_if_if_for_equal_tmp_5_1 | while_else_4_if_if_for_equal_tmp_6_1
      | while_else_4_if_if_for_equal_tmp_7_1 | and_515_cse | while_else_4_if_if_for_equal_tmp_9_1
      | while_else_4_if_if_for_equal_tmp_10_1 | while_else_4_if_if_for_equal_tmp_11_1
      | while_else_4_if_if_for_equal_tmp_12_1 | while_else_4_if_if_for_equal_tmp_13_1
      | while_else_4_if_if_for_while_else_4_if_if_for_and_13_itm_1 | while_else_4_if_if_for_while_else_4_if_if_for_and_14_itm_1))
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_or_16_cse_1 = if_axi_rd_ar_PopNB_mioi_bawt | (~((~ while_asn_25_itm_1)
      & while_stage_v_1));
  assign while_or_17_cse_1 = if_axi_wr_aw_PopNB_mioi_bawt | (~((~ while_asn_30_itm_1)
      & while_stage_v_1));
  assign while_or_18_cse_1 = regIn_PopNB_mioi_bawt | (~((~ while_asn_34_itm_1) &
      while_stage_v_1));
  assign while_or_19_cse_1 = if_axi_wr_w_PopNB_mioi_bawt | (~(operator_3_false_2_operator_3_false_2_and_svs_st_1
      & (~ operator_3_false_1_operator_3_false_1_and_svs_st_1) & while_stage_v_1));
  assign while_nand_2_cse = ~(operator_3_false_1_operator_3_false_1_and_svs_st_2
      & while_stage_v_2);
  assign while_or_cse_1 = if_axi_rd_r_Push_mioi_bawt | while_nand_2_cse;
  assign while_or_14_cse_1 = if_axi_wr_b_Push_mioi_bawt | (~(while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
      & operator_3_false_2_operator_3_false_2_and_svs_st_2 & (~ operator_3_false_1_operator_3_false_1_and_svs_st_2)
      & while_stage_v_2));
  assign while_else_4_if_if_if_1_old_data_sva_1 = MUX_v_64_14_2(reg_0_sva_mx1, reg_1_sva_mx1,
      reg_2_sva_mx1, reg_3_sva_mx1, reg_4_sva_mx1, reg_5_sva_mx1, reg_6_sva_mx1,
      reg_7_sva_mx1, reg_8_sva_mx1, reg_9_sva_mx1, reg_10_sva_mx1, reg_11_sva_mx1,
      reg_12_sva_mx1, reg_13_sva_mx1, while_else_4_if_if_regAddr_acc_itm_6_3);
  assign arb_pick_if_1_not_15 = nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm_mx0w0
      & (~(arb_pick_priority_4_sva_mx0w0 | nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm_mx0w0));
  assign while_and_31_nl = if_axi_rd_ar_PopNB_mioi_ivld_mxwt & (~ read_arb_req_sva);
  assign while_mux_17_tmp = MUX_v_8_2_2(axiRdLen_sva, (if_axi_rd_ar_PopNB_mioi_idat_mxwt[27:20]),
      while_and_31_nl);
  assign while_mux_32_tmp = MUX_v_4_2_2((regIn_PopNB_mioi_idat_mxwt[3:0]), regwr_addr_6_3_sva,
      regIn_arb_req_sva);
  assign and_dcpl = operator_3_false_1_operator_3_false_1_and_svs_st_1 & while_stage_v_1;
  assign or_dcpl_2 = regIn_PopNB_mioi_bawt | while_asn_34_itm_1;
  assign or_dcpl_3 = if_axi_wr_aw_PopNB_mioi_bawt | while_asn_30_itm_1;
  assign or_dcpl_4 = if_axi_rd_ar_PopNB_mioi_bawt | while_asn_25_itm_1;
  assign mux_5_cse = MUX_s_1_2_2(nand_142_cse_1, if_axi_rd_r_Push_mioi_bawt, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign or_tmp_54 = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_9_1) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign or_68_cse = (~ (regwr_addr_6_3_sva[3])) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | operator_3_false_1_operator_3_false_1_and_svs_2 | mux_5_cse;
  assign mux_83_nl = MUX_s_1_2_2(or_68_cse, or_tmp_54, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_10 = ~(while_stage_v_2 & (~ mux_83_nl));
  assign nor_70_cse = ~((~ (regwr_addr_6_3_sva[3])) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | operator_3_false_1_operator_3_false_1_and_svs_2);
  assign or_662_cse = nor_70_cse | mux_5_cse;
  assign mux_tmp_86 = MUX_s_1_2_2(or_662_cse, (~ or_tmp_54), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_tmp_87 = MUX_s_1_2_2((~ mux_tmp_86), nand_tmp_10, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign or_661_nl = (~((~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_9_1) | operator_3_false_1_operator_3_false_1_and_svs_2))
      | mux_5_cse;
  assign mux_88_nl = MUX_s_1_2_2(or_662_cse, or_661_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_14 = ~(while_stage_v_2 & (~ mux_88_nl));
  assign or_tmp_70 = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_10_1) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign mux_109_nl = MUX_s_1_2_2(or_68_cse, or_tmp_70, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_15 = ~(while_stage_v_2 & (~ mux_109_nl));
  assign mux_tmp_112 = MUX_s_1_2_2(or_662_cse, (~ or_tmp_70), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nor_136_cse = ~(nor_70_cse | mux_5_cse);
  assign nor_137_nl = ~((~((~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_10_1) | operator_3_false_1_operator_3_false_1_and_svs_2))
      | mux_5_cse);
  assign mux_114_nl = MUX_s_1_2_2(nor_136_cse, nor_137_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_19 = ~(while_stage_v_2 & mux_114_nl);
  assign or_tmp_86 = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_6_1) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign or_100_cse = (regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (~ (regwr_addr_6_3_sva[2])) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign mux_133_nl = MUX_s_1_2_2(or_100_cse, or_tmp_86, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_20 = ~(while_stage_v_2 & (~ mux_133_nl));
  assign or_668_cse = nor_97_cse | mux_5_cse;
  assign mux_tmp_136 = MUX_s_1_2_2(or_668_cse, (~ or_tmp_86), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_302_cse = operator_3_false_2_operator_3_false_2_and_svs_st_2 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
      & while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1 & (~ if_axi_wr_b_Push_mioi_bawt);
  assign or_113_nl = and_302_cse | (~ operator_3_false_3_operator_3_false_3_and_svs_1)
      | (while_mux_32_tmp[3:2]!=2'b01);
  assign nand_128_nl = ~(if_axi_rd_r_Push_mioi_bawt & operator_3_false_3_operator_3_false_3_and_svs_1
      & (while_mux_32_tmp[3:2]==2'b01));
  assign mux_tmp_143 = MUX_s_1_2_2(or_113_nl, nand_128_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign or_tmp_103 = (~ operator_3_false_3_operator_3_false_3_and_svs_1) | (while_mux_32_tmp[3:2]!=2'b01);
  assign and_14_nl = nand_142_cse_1 & or_tmp_103;
  assign and_13_nl = if_axi_rd_r_Push_mioi_bawt & or_tmp_103;
  assign mux_tmp_144 = MUX_s_1_2_2(and_14_nl, and_13_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_148_nl = MUX_s_1_2_2(mux_151_cse, or_tmp_86, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_tmp_149 = MUX_s_1_2_2(or_tmp_103, mux_148_nl, while_stage_v_2);
  assign or_tmp_114 = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_11_1) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign mux_165_nl = MUX_s_1_2_2(or_68_cse, or_tmp_114, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_26 = ~(while_stage_v_2 & (~ mux_165_nl));
  assign mux_tmp_168 = MUX_s_1_2_2(or_662_cse, (~ or_tmp_114), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_tmp_169 = MUX_s_1_2_2((~ mux_tmp_168), nand_tmp_26, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign nor_139_nl = ~((~((~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_11_1) | operator_3_false_1_operator_3_false_1_and_svs_2))
      | mux_5_cse);
  assign mux_170_nl = MUX_s_1_2_2(nor_136_cse, nor_139_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_30 = ~(while_stage_v_2 & mux_170_nl);
  assign or_tmp_129 = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_3_1) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign or_143_cse = (regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | operator_3_false_1_operator_3_false_1_and_svs_2 | mux_5_cse;
  assign mux_191_nl = MUX_s_1_2_2(or_143_cse, or_tmp_129, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_31 = ~(while_stage_v_2 & (~ mux_191_nl));
  assign nor_81_cse = ~((regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | operator_3_false_1_operator_3_false_1_and_svs_2);
  assign or_673_cse = nor_81_cse | mux_5_cse;
  assign mux_tmp_194 = MUX_s_1_2_2(or_673_cse, (~ or_tmp_129), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_tmp_195 = MUX_s_1_2_2((~ mux_tmp_194), nand_tmp_31, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign or_672_nl = (~((~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_3_1) | operator_3_false_1_operator_3_false_1_and_svs_2))
      | mux_5_cse;
  assign mux_196_nl = MUX_s_1_2_2(or_673_cse, or_672_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_35 = ~(while_stage_v_2 & (~ mux_196_nl));
  assign or_tmp_145 = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_7_1) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign mux_217_nl = MUX_s_1_2_2(or_100_cse, or_tmp_145, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_36 = ~(while_stage_v_2 & (~ mux_217_nl));
  assign mux_tmp_220 = MUX_s_1_2_2(or_668_cse, (~ or_tmp_145), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_tmp_221 = MUX_s_1_2_2((~ mux_tmp_220), nand_tmp_36, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_233_nl = MUX_s_1_2_2(mux_151_cse, or_tmp_145, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_tmp_234 = MUX_s_1_2_2(or_tmp_103, mux_233_nl, while_stage_v_2);
  assign or_tmp_172 = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_12_1) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign mux_250_nl = MUX_s_1_2_2(or_68_cse, or_tmp_172, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_42 = ~(while_stage_v_2 & (~ mux_250_nl));
  assign mux_tmp_253 = MUX_s_1_2_2(or_662_cse, (~ or_tmp_172), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nor_141_nl = ~((~((~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_12_1) | operator_3_false_1_operator_3_false_1_and_svs_2))
      | mux_5_cse);
  assign mux_255_nl = MUX_s_1_2_2(nor_136_cse, nor_141_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_46 = ~(while_stage_v_2 & mux_255_nl);
  assign or_tmp_188 = (~ while_else_4_if_if_for_equal_tmp_13_1) | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | operator_3_false_1_operator_3_false_1_and_svs_2 | mux_5_cse;
  assign mux_274_nl = MUX_s_1_2_2(or_68_cse, or_tmp_188, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_47 = ~(while_stage_v_2 & (~ mux_274_nl));
  assign mux_tmp_277 = MUX_s_1_2_2(or_662_cse, (~ or_tmp_188), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_tmp_278 = MUX_s_1_2_2((~ mux_tmp_277), nand_tmp_47, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign nor_143_nl = ~((~((~ while_else_4_if_if_for_equal_tmp_13_1) | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | operator_3_false_1_operator_3_false_1_and_svs_2)) | mux_5_cse);
  assign mux_279_nl = MUX_s_1_2_2(nor_136_cse, nor_143_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_51 = ~(while_stage_v_2 & mux_279_nl);
  assign or_tmp_204 = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_5_1) | operator_3_false_1_operator_3_false_1_and_svs_2
      | mux_5_cse;
  assign mux_300_nl = MUX_s_1_2_2(or_143_cse, or_tmp_204, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_52 = ~(while_stage_v_2 & (~ mux_300_nl));
  assign mux_tmp_303 = MUX_s_1_2_2(or_673_cse, (~ or_tmp_204), operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_tmp_304 = MUX_s_1_2_2((~ mux_tmp_303), nand_tmp_52, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign nor_144_nl = ~(nor_81_cse | mux_5_cse);
  assign nor_145_nl = ~((~((~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_5_1) | operator_3_false_1_operator_3_false_1_and_svs_2))
      | mux_5_cse);
  assign mux_305_nl = MUX_s_1_2_2(nor_144_nl, nor_145_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nand_tmp_56 = ~(while_stage_v_2 & mux_305_nl);
  assign or_235_nl = if_axi_wr_b_Push_mioi_bawt | nand_198_cse;
  assign mux_325_nl = MUX_s_1_2_2(or_235_nl, if_axi_rd_r_Push_mioi_bawt, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign or_dcpl_17 = mux_325_nl | (~ while_stage_v_2);
  assign or_234_cse = if_axi_wr_w_PopNB_mioi_bawt | (~ operator_3_false_2_operator_3_false_2_and_svs_st_1)
      | operator_3_false_1_operator_3_false_1_and_svs_st_1;
  assign or_tmp_221 = (~ operator_3_false_2_operator_3_false_2_and_svs_st_2) | (~
      while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1)
      | (~ while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1) | if_axi_wr_b_Push_mioi_bawt
      | operator_3_false_1_operator_3_false_1_and_svs_st_2 | (~ while_stage_v_2);
  assign and_305_cse = operator_3_false_2_operator_3_false_2_and_svs_st_1 & if_axi_wr_w_PopNB_mioi_ivld_mxwt
      & if_axi_wr_w_PopNB_mioi_bawt;
  assign or_tmp_228 = (~ while_stage_v_2) | operator_3_false_1_operator_3_false_1_and_svs_st_2
      | operator_3_false_1_operator_3_false_1_and_svs_2 | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ operator_3_false_2_operator_3_false_2_and_svs_2) | while_else_4_if_if_while_else_4_if_if_nand_tmp_1
      | (~ operator_3_false_2_operator_3_false_2_and_svs_st_2) | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1)
      | (~ while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1) | if_axi_wr_b_Push_mioi_bawt;
  assign or_tmp_234 = (~ while_stage_v_2) | operator_3_false_1_operator_3_false_1_and_svs_st_2
      | operator_3_false_1_operator_3_false_1_and_svs_2 | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ operator_3_false_2_operator_3_false_2_and_svs_2) | (~ operator_3_false_2_operator_3_false_2_and_svs_st_2)
      | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1)
      | (~ while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1) | if_axi_wr_b_Push_mioi_bawt;
  assign and_dcpl_19 = operator_3_false_2_operator_3_false_2_and_svs_st_1 & (~ operator_3_false_1_operator_3_false_1_and_svs_st_1)
      & while_stage_v_1;
  assign and_dcpl_20 = (if_axi_wr_w_PopNB_mioi_idat_mxwt[64]) & if_axi_wr_w_PopNB_mioi_bawt;
  assign nor_tmp_25 = while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
      & operator_3_false_2_operator_3_false_2_and_svs_st_2;
  assign or_293_nl = if_axi_wr_b_Push_mioi_bawt | (~ nor_tmp_25);
  assign mux_tmp_364 = MUX_s_1_2_2(or_293_nl, if_axi_rd_r_Push_mioi_bawt, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign or_dcpl_25 = mux_tmp_364 | (~ while_stage_v_2);
  assign and_dcpl_24 = or_dcpl_25 & or_dcpl_4;
  assign and_dcpl_25 = and_dcpl_24 & or_dcpl_3;
  assign and_dcpl_26 = and_dcpl_25 & or_dcpl_2;
  assign or_dcpl_28 = (~(if_axi_wr_w_PopNB_mioi_bawt & operator_3_false_2_operator_3_false_2_and_svs_st_1))
      | operator_3_false_1_operator_3_false_1_and_svs_st_1 | (~ while_stage_v_1);
  assign and_dcpl_32 = ~(regIn_PopNB_mioi_bawt | while_asn_34_itm_1);
  assign and_dcpl_33 = ~(if_axi_wr_aw_PopNB_mioi_bawt | while_asn_30_itm_1);
  assign and_dcpl_34 = ~(if_axi_rd_ar_PopNB_mioi_bawt | while_asn_25_itm_1);
  assign and_dcpl_35 = (~ mux_tmp_364) & while_stage_v_2;
  assign or_dcpl_35 = ~(operator_3_false_1_operator_3_false_1_and_svs_st_1 & while_stage_v_1);
  assign or_dcpl_36 = and_dcpl_33 | and_dcpl_32;
  assign or_dcpl_38 = and_dcpl_35 | and_dcpl_34;
  assign or_dcpl_39 = or_dcpl_38 | or_dcpl_36 | or_dcpl_35;
  assign or_tmp_280 = select_mask_0_sva | (~ select_mask_2_1_sva_0) | select_mask_2_1_sva_1;
  assign or_tmp_282 = (~ if_axi_wr_aw_PopNB_mioi_ivld_mxwt) | while_asn_30_itm_1;
  assign not_tmp_228 = ~(if_axi_wr_aw_PopNB_mioi_bawt & and_dcpl_24);
  assign nor_106_nl = ~(or_tmp_282 | not_tmp_228);
  assign mux_tmp_370 = MUX_s_1_2_2(nor_106_nl, and_dcpl_25, write_arb_req_sva);
  assign and_tmp_19 = or_dcpl_2 & mux_tmp_370;
  assign and_73_nl = while_asn_34_itm_1 & mux_tmp_370;
  assign mux_371_nl = MUX_s_1_2_2(and_tmp_19, and_73_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign or_tmp_285 = regIn_arb_req_sva | (~ mux_371_nl);
  assign or_tmp_287 = read_arb_req_sva | and_dcpl_35;
  assign or_330_nl = while_while_or_tmp | (~(if_axi_rd_ar_PopNB_mioi_bawt & or_dcpl_25));
  assign mux_tmp_373 = MUX_s_1_2_2(or_330_nl, or_tmp_287, while_asn_25_itm_1);
  assign nand_tmp_63 = ~(or_dcpl_3 & (~ mux_tmp_373));
  assign or_690_nl = (~ if_axi_wr_aw_PopNB_mioi_ivld_mxwt) | while_asn_30_itm_1 |
      (~ if_axi_wr_aw_PopNB_mioi_bawt) | mux_tmp_373;
  assign mux_374_itm = MUX_s_1_2_2(or_690_nl, nand_tmp_63, write_arb_req_sva);
  assign nand_tmp_66 = ~(or_dcpl_2 & (~ mux_374_itm));
  assign or_322_nl = or_tmp_280 | (~ and_dcpl_26);
  assign nand_65_nl = ~(while_asn_34_itm_1 & (~ mux_374_itm));
  assign mux_375_nl = MUX_s_1_2_2(nand_tmp_66, nand_65_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign or_332_nl = regIn_arb_req_sva | mux_375_nl;
  assign mux_372_nl = MUX_s_1_2_2((~ and_tmp_19), or_tmp_285, arb_next_1_2_sva);
  assign mux_376_nl = MUX_s_1_2_2(or_332_nl, mux_372_nl, arb_next_1_1_sva);
  assign mux_tmp_378 = MUX_s_1_2_2(or_322_nl, mux_376_nl, arb_needs_update_sva);
  assign or_tmp_292 = (~ arb_next_1_1_sva) | arb_next_1_2_sva;
  assign mux_tmp_381 = MUX_s_1_2_2((~ and_tmp_19), or_tmp_285, or_tmp_292);
  assign nor_tmp_28 = ~(operator_3_false_1_operator_3_false_1_and_svs_st_1 | (~ operator_3_false_2_operator_3_false_2_and_svs_st_1));
  assign nor_tmp_30 = arb_next_1_2_sva & regIn_arb_req_sva;
  assign and_dcpl_55 = (~ operator_3_false_1_operator_3_false_1_and_svs_st_1) & while_stage_v_1;
  assign and_dcpl_58 = and_dcpl_26 & if_axi_wr_w_PopNB_mioi_bawt & operator_3_false_2_operator_3_false_2_and_svs_st_1
      & and_dcpl_55;
  assign nand_tmp_71 = ~(while_stage_v_2 & (~ mux_5_cse));
  assign and_tmp_21 = or_dcpl_3 & nand_tmp_71;
  assign or_351_nl = regIn_PopNB_mioi_ivld_mxwt | (~(regIn_PopNB_mioi_bawt & and_tmp_21));
  assign mux_398_nl = MUX_s_1_2_2(or_351_nl, (~ and_tmp_21), while_asn_34_itm_1);
  assign or_tmp_311 = regIn_arb_req_sva | mux_398_nl;
  assign or_tmp_315 = while_stage_v_1 | regIn_arb_req_sva | (~ nand_tmp_71);
  assign and_68_nl = while_asn_30_itm_1 & and_dcpl_24;
  assign mux_404_itm = MUX_s_1_2_2(and_dcpl_25, and_68_nl, if_axi_wr_aw_PopNB_mioi_ivld_mxwt);
  assign or_tmp_322 = (~ or_dcpl_2) | write_arb_req_sva | (~ mux_404_itm);
  assign and_tmp_26 = or_dcpl_2 & or_dcpl_3 & nand_tmp_71;
  assign and_333_nl = operator_8_false_operator_8_false_nor_mdf_sva & or_28_cse &
      and_tmp_26;
  assign nor_107_nl = ~((while_mux_17_tmp!=8'b00000000) | (~ and_tmp_26));
  assign mux_413_nl = MUX_s_1_2_2(and_333_nl, nor_107_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign nand_tmp_74 = ~(operator_3_false_1_operator_3_false_1_and_svs_1 & mux_413_nl);
  assign not_tmp_258 = ~(or_234_cse & and_tmp_26);
  assign or_dcpl_43 = ~(mux_tmp_364 & while_stage_v_2);
  assign nand_78_nl = ~(while_asn_30_itm_1 & (~ mux_tmp_373));
  assign mux_tmp_423 = MUX_s_1_2_2(nand_tmp_63, nand_78_nl, if_axi_wr_aw_PopNB_mioi_ivld_mxwt);
  assign and_tmp_32 = read_arb_req_sva & or_dcpl_25;
  assign and_107_nl = while_while_or_tmp & if_axi_rd_ar_PopNB_mioi_bawt & or_dcpl_25;
  assign mux_tmp_424 = MUX_s_1_2_2(and_107_nl, and_tmp_32, while_asn_25_itm_1);
  assign and_tmp_33 = or_dcpl_3 & mux_tmp_424;
  assign and_335_nl = if_axi_wr_aw_PopNB_mioi_bawt & (~ mux_tmp_373);
  assign mux_425_nl = MUX_s_1_2_2(and_335_nl, mux_tmp_424, while_asn_30_itm_1);
  assign mux_426_nl = MUX_s_1_2_2(and_tmp_33, mux_425_nl, if_axi_wr_aw_PopNB_mioi_ivld_mxwt);
  assign mux_tmp_427 = MUX_s_1_2_2((~ mux_426_nl), nand_tmp_63, write_arb_req_sva);
  assign or_tmp_349 = (~ regIn_PopNB_mioi_bawt) | write_arb_req_sva;
  assign nand_tmp_80 = ~(or_dcpl_2 & (~ mux_tmp_427));
  assign or_394_nl = or_tmp_349 | mux_tmp_423;
  assign mux_428_nl = MUX_s_1_2_2(or_394_nl, mux_tmp_427, while_asn_34_itm_1);
  assign mux_429_nl = MUX_s_1_2_2(nand_tmp_80, mux_428_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign or_391_nl = (~ or_dcpl_2) | write_arb_req_sva | mux_tmp_423;
  assign mux_430_nl = MUX_s_1_2_2(mux_429_nl, or_391_nl, regIn_arb_req_sva);
  assign mux_tmp_431 = ~(arb_needs_update_sva & (~ mux_430_nl));
  assign nor_110_nl = ~(or_tmp_349 | (~ mux_404_itm));
  assign mux_434_nl = MUX_s_1_2_2(nor_110_nl, mux_tmp_370, while_asn_34_itm_1);
  assign mux_435_nl = MUX_s_1_2_2(and_tmp_19, mux_434_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign mux_tmp_437 = MUX_s_1_2_2((~ mux_435_nl), or_tmp_322, regIn_arb_req_sva);
  assign nand_tmp_85 = ~(or_dcpl_2 & (~ nand_tmp_63));
  assign and_tmp_36 = or_dcpl_2 & and_tmp_33;
  assign mux_957_nl = MUX_s_1_2_2(mux_tmp_431, nand_tmp_80, operator_3_false_3_operator_3_false_3_and_svs_1);
  assign mux_453_nl = MUX_s_1_2_2(mux_957_nl, mux_tmp_431, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_685_nl = MUX_s_1_2_2(mux_tmp_431, nand_tmp_80, operator_3_false_3_operator_3_false_3_and_svs_1);
  assign and_337_nl = regIn_PopNB_mioi_bawt & (~ nand_tmp_63);
  assign mux_443_nl = MUX_s_1_2_2(and_337_nl, and_tmp_33, while_asn_34_itm_1);
  assign mux_444_nl = MUX_s_1_2_2(and_tmp_36, mux_443_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign mux_445_nl = MUX_s_1_2_2((~ mux_444_nl), nand_tmp_85, regIn_arb_req_sva);
  assign mux_447_nl = MUX_s_1_2_2(mux_tmp_431, mux_445_nl, and_352_cse);
  assign mux_450_nl = MUX_s_1_2_2(mux_685_nl, mux_447_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nand_88_nl = ~(if_axi_wr_w_PopNB_mioi_bawt & (~ mux_450_nl));
  assign mux_454_nl = MUX_s_1_2_2(mux_453_nl, nand_88_nl, nor_tmp_28);
  assign nand_83_nl = ~(or_28_cse & (~ mux_tmp_431));
  assign nand_82_nl = ~(or_28_cse & (~ mux_tmp_437));
  assign mux_439_nl = MUX_s_1_2_2(nand_83_nl, nand_82_nl, operator_8_false_operator_8_false_nor_mdf_sva);
  assign mux_438_nl = MUX_s_1_2_2(mux_tmp_437, mux_tmp_431, or_310_cse);
  assign mux_440_nl = MUX_s_1_2_2(mux_439_nl, mux_438_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_tmp_455 = MUX_s_1_2_2(mux_454_nl, mux_440_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign or_tmp_368 = (~ while_asn_34_itm_1) | write_arb_req_sva;
  assign or_tmp_369 = ~(while_asn_30_itm_1 | (~ if_axi_wr_aw_PopNB_mioi_ivld_mxwt));
  assign or_tmp_370 = (~(while_asn_25_itm_1 | (~ if_axi_rd_ar_PopNB_mioi_ivld_mxwt)))
      | read_arb_req_sva;
  assign or_tmp_371 = or_tmp_369 | or_tmp_370;
  assign or_421_nl = if_axi_wr_aw_PopNB_mioi_ivld_mxwt | or_tmp_370;
  assign mux_460_nl = MUX_s_1_2_2(or_421_nl, or_tmp_370, while_asn_30_itm_1);
  assign or_tmp_377 = write_arb_req_sva | mux_460_nl;
  assign or_418_nl = write_arb_req_sva | or_tmp_371;
  assign mux_461_nl = MUX_s_1_2_2(or_tmp_377, or_418_nl, while_asn_34_itm_1);
  assign or_417_nl = or_tmp_368 | or_tmp_371;
  assign mux_462_nl = MUX_s_1_2_2(mux_461_nl, or_417_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign or_tmp_378 = regIn_arb_req_sva | mux_462_nl;
  assign or_427_nl = write_arb_req_sva | or_tmp_369;
  assign mux_464_nl = MUX_s_1_2_2(while_while_or_1_tmp, or_427_nl, while_asn_34_itm_1);
  assign or_426_nl = or_tmp_368 | or_tmp_369;
  assign mux_465_nl = MUX_s_1_2_2(mux_464_nl, or_426_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign or_tmp_384 = regIn_arb_req_sva | mux_465_nl;
  assign or_tmp_385 = (~ operator_3_false_2_operator_3_false_2_and_svs_st_1) | operator_3_false_1_operator_3_false_1_and_svs_st_1;
  assign or_436_nl = regIn_arb_req_sva | write_arb_req_sva | read_arb_req_sva;
  assign mux_478_nl = MUX_s_1_2_2(or_tmp_378, or_tmp_377, operator_3_false_3_operator_3_false_3_and_svs_1);
  assign or_434_nl = (~ while_asn_34_itm_1) | or_tmp_370;
  assign mux_475_nl = MUX_s_1_2_2(or_tmp_370, or_434_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign or_435_nl = regIn_arb_req_sva | mux_475_nl;
  assign mux_476_nl = MUX_s_1_2_2(or_tmp_378, or_435_nl, and_352_cse);
  assign mux_477_nl = MUX_s_1_2_2(mux_476_nl, or_tmp_378, or_tmp_385);
  assign mux_479_nl = MUX_s_1_2_2(mux_478_nl, mux_477_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_467_nl = MUX_s_1_2_2(or_tmp_378, or_tmp_384, operator_8_false_operator_8_false_nor_mdf_sva);
  assign mux_466_nl = MUX_s_1_2_2(or_tmp_384, or_tmp_378, or_310_cse);
  assign mux_468_nl = MUX_s_1_2_2(mux_467_nl, mux_466_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_480_nl = MUX_s_1_2_2(mux_479_nl, mux_468_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign mux_481_itm = MUX_s_1_2_2(or_436_nl, mux_480_nl, while_stage_v_1);
  assign and_dcpl_77 = operator_3_false_1_operator_3_false_1_and_svs_1 & while_stage_v_1;
  assign and_dcpl_78 = and_dcpl_26 & or_234_cse;
  assign and_dcpl_79 = and_dcpl_78 & and_dcpl_77;
  assign and_dcpl_80 = (~ operator_3_false_1_operator_3_false_1_and_svs_1) & while_stage_v_1;
  assign and_dcpl_81 = and_dcpl_78 & and_dcpl_80;
  assign and_dcpl_83 = (~ if_axi_wr_w_PopNB_mioi_bawt) & operator_3_false_2_operator_3_false_2_and_svs_st_1
      & (~ operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign and_tmp_39 = or_dcpl_3 & or_dcpl_4 & or_dcpl_2 & nand_tmp_71;
  assign and_tmp_40 = or_234_cse & and_tmp_39;
  assign and_130_nl = arb_needs_update_sva & nand_tmp_71;
  assign and_129_nl = operator_3_false_3_operator_3_false_3_and_svs_1 & and_tmp_40;
  assign and_127_nl = (if_axi_wr_w_PopNB_mioi_idat_mxwt[64]) & if_axi_wr_w_PopNB_mioi_ivld_mxwt
      & if_axi_wr_w_PopNB_mioi_bawt & and_tmp_39;
  assign mux_484_nl = MUX_s_1_2_2(and_tmp_39, and_127_nl, nor_tmp_28);
  assign mux_485_nl = MUX_s_1_2_2(and_129_nl, mux_484_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign and_341_nl = operator_8_false_operator_8_false_nor_mdf_sva & or_28_cse &
      and_tmp_39;
  assign nor_111_nl = ~((while_mux_17_tmp!=8'b00000000) | (~ and_tmp_39));
  assign mux_483_nl = MUX_s_1_2_2(and_341_nl, nor_111_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_486_nl = MUX_s_1_2_2(mux_485_nl, mux_483_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign mux_487_nl = MUX_s_1_2_2(mux_486_nl, and_tmp_40, arb_needs_update_sva);
  assign mux_488_itm = MUX_s_1_2_2(and_130_nl, mux_487_nl, while_stage_v_1);
  assign mux_489_itm = MUX_s_1_2_2(or_dcpl_25, and_dcpl_78, while_stage_v_1);
  assign or_dcpl_51 = while_asn_25_itm_1 | (~ if_axi_rd_ar_PopNB_mioi_ivld_mxwt)
      | read_arb_req_sva;
  assign and_343_nl = or_28_cse & ((~ operator_3_false_1_operator_3_false_1_and_svs_1)
      | operator_8_false_operator_8_false_nor_mdf_sva) & nand_tmp_71;
  assign nor_114_nl = ~((while_mux_17_tmp!=8'b00000000) | (~ nand_tmp_71));
  assign mux_496_nl = MUX_s_1_2_2(nand_tmp_71, nor_114_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign mux_497_nl = MUX_s_1_2_2(and_343_nl, mux_496_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign and_dcpl_91 = mux_497_nl & or_dcpl_4 & or_dcpl_3 & or_dcpl_2 & while_stage_v_1;
  assign or_dcpl_52 = or_tmp_282 | write_arb_req_sva;
  assign or_tmp_435 = (~ select_mask_0_sva) | select_mask_2_1_sva_0 | select_mask_2_1_sva_1;
  assign mux_517_nl = MUX_s_1_2_2(not_tmp_228, mux_tmp_373, while_asn_30_itm_1);
  assign mux_518_nl = MUX_s_1_2_2(nand_tmp_63, mux_517_nl, if_axi_wr_aw_PopNB_mioi_ivld_mxwt);
  assign mux_tmp_519 = MUX_s_1_2_2((~ mux_518_nl), and_dcpl_25, write_arb_req_sva);
  assign and_tmp_60 = regIn_PopNB_mioi_bawt & and_dcpl_25;
  assign and_tmp_61 = or_dcpl_2 & mux_tmp_519;
  assign mux_524_nl = MUX_s_1_2_2((~ and_tmp_60), nand_tmp_63, while_asn_34_itm_1);
  assign mux_525_nl = MUX_s_1_2_2(nand_tmp_85, mux_524_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign mux_526_nl = MUX_s_1_2_2((~ mux_525_nl), and_dcpl_26, regIn_arb_req_sva);
  assign mux_tmp_527 = MUX_s_1_2_2((~ nand_tmp_85), mux_526_nl, arb_next_1_2_sva);
  assign and_161_nl = or_tmp_435 & and_dcpl_26;
  assign mux_520_nl = MUX_s_1_2_2(and_tmp_60, mux_tmp_519, while_asn_34_itm_1);
  assign mux_521_nl = MUX_s_1_2_2(and_tmp_61, mux_520_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign mux_522_nl = MUX_s_1_2_2(mux_521_nl, and_dcpl_26, regIn_arb_req_sva);
  assign mux_523_nl = MUX_s_1_2_2(and_tmp_61, mux_522_nl, arb_next_1_2_sva);
  assign mux_528_nl = MUX_s_1_2_2(mux_tmp_527, mux_523_nl, arb_next_1_1_sva);
  assign mux_tmp_530 = MUX_s_1_2_2(and_161_nl, mux_528_nl, arb_needs_update_sva);
  assign mux_537_nl = MUX_s_1_2_2((~ nand_tmp_85), and_tmp_61, arb_next_1_1_sva);
  assign mux_683_itm = MUX_s_1_2_2(mux_tmp_530, mux_537_nl, operator_3_false_3_operator_3_false_3_and_svs_1);
  assign mux_543_nl = MUX_s_1_2_2(mux_683_itm, mux_tmp_530, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_535_nl = MUX_s_1_2_2(mux_tmp_530, mux_tmp_527, and_352_cse);
  assign mux_540_nl = MUX_s_1_2_2(mux_683_itm, mux_535_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign and_166_nl = if_axi_wr_w_PopNB_mioi_bawt & mux_540_nl;
  assign mux_544_nl = MUX_s_1_2_2(mux_543_nl, and_166_nl, nor_tmp_28);
  assign and_165_nl = or_28_cse & mux_tmp_530;
  assign and_164_nl = or_28_cse & and_dcpl_26;
  assign mux_532_nl = MUX_s_1_2_2(and_165_nl, and_164_nl, operator_8_false_operator_8_false_nor_mdf_sva);
  assign mux_531_nl = MUX_s_1_2_2(and_dcpl_26, mux_tmp_530, or_310_cse);
  assign mux_533_nl = MUX_s_1_2_2(mux_532_nl, mux_531_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_tmp_545 = MUX_s_1_2_2(mux_544_nl, mux_533_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign or_tmp_439 = nor_tmp_30 | write_arb_req_sva;
  assign and_170_nl = while_asn_30_itm_1 & mux_tmp_424;
  assign mux_555_itm = MUX_s_1_2_2(and_tmp_33, and_170_nl, if_axi_wr_aw_PopNB_mioi_ivld_mxwt);
  assign or_tmp_456 = (~ or_dcpl_2) | write_arb_req_sva | (~ mux_555_itm);
  assign and_171_nl = while_asn_34_itm_1 & and_tmp_33;
  assign mux_558_nl = MUX_s_1_2_2(and_tmp_36, and_171_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign or_520_nl = regIn_arb_req_sva | (~ mux_558_nl);
  assign mux_tmp_559 = MUX_s_1_2_2((~ and_tmp_36), or_520_nl, arb_next_1_2_sva);
  assign or_513_nl = or_tmp_435 | (~ and_dcpl_26);
  assign or_515_nl = or_tmp_368 | (~ mux_555_itm);
  assign mux_556_nl = MUX_s_1_2_2(or_tmp_456, or_515_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign or_519_nl = regIn_arb_req_sva | mux_556_nl;
  assign mux_557_nl = MUX_s_1_2_2(or_tmp_456, or_519_nl, arb_next_1_2_sva);
  assign mux_560_nl = MUX_s_1_2_2(mux_tmp_559, mux_557_nl, arb_next_1_1_sva);
  assign mux_tmp_562 = MUX_s_1_2_2(or_513_nl, mux_560_nl, arb_needs_update_sva);
  assign nor_116_cse = ~((while_mux_17_tmp!=8'b00000000));
  assign mux_567_nl = MUX_s_1_2_2((~ and_tmp_36), or_tmp_456, arb_next_1_1_sva);
  assign mux_684_itm = MUX_s_1_2_2(mux_tmp_562, mux_567_nl, operator_3_false_3_operator_3_false_3_and_svs_1);
  assign mux_573_nl = MUX_s_1_2_2(mux_684_itm, mux_tmp_562, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_565_nl = MUX_s_1_2_2(mux_tmp_562, mux_tmp_559, and_352_cse);
  assign mux_570_nl = MUX_s_1_2_2(mux_684_itm, mux_565_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nand_97_nl = ~(if_axi_wr_w_PopNB_mioi_bawt & (~ mux_570_nl));
  assign mux_574_nl = MUX_s_1_2_2(mux_573_nl, nand_97_nl, nor_tmp_28);
  assign or_522_nl = operator_8_false_operator_8_false_nor_mdf_sva | (~(or_28_cse
      & (~ mux_tmp_562)));
  assign or_692_nl = nor_116_cse | mux_tmp_562;
  assign mux_563_nl = MUX_s_1_2_2(or_522_nl, or_692_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_tmp_575 = MUX_s_1_2_2(mux_574_nl, mux_563_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign and_dcpl_117 = nor_tmp_25 & while_stage_v_2 & (~ if_axi_wr_b_Push_mioi_bawt)
      & (~ operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign or_dcpl_64 = (~ nor_tmp_25) | (~ while_stage_v_2) | if_axi_wr_b_Push_mioi_bawt
      | operator_3_false_1_operator_3_false_1_and_svs_st_2;
  assign nand_tmp_98 = ~(while_stage_v_2 & (~ mux_tmp_364));
  assign and_tmp_70 = or_dcpl_4 & nand_tmp_98;
  assign and_tmp_71 = if_axi_wr_aw_PopNB_mioi_bawt & and_tmp_70;
  assign and_tmp_72 = or_dcpl_3 & and_tmp_70;
  assign and_tmp_75 = regIn_PopNB_mioi_bawt & and_tmp_72;
  assign and_tmp_76 = or_dcpl_2 & and_tmp_72;
  assign nor_119_nl = ~(if_axi_wr_aw_PopNB_mioi_ivld_mxwt | (~ and_tmp_71));
  assign mux_610_itm = MUX_s_1_2_2(nor_119_nl, and_tmp_70, while_asn_30_itm_1);
  assign or_tmp_509 = (~ or_dcpl_2) | write_arb_req_sva | (~ mux_610_itm);
  assign or_tmp_510 = read_arb_req_sva | (~ nand_tmp_98);
  assign or_581_nl = (~ if_axi_rd_ar_PopNB_mioi_bawt) | if_axi_rd_ar_PopNB_mioi_ivld_mxwt
      | read_arb_req_sva | (~ nand_tmp_98);
  assign mux_tmp_611 = MUX_s_1_2_2(or_581_nl, or_tmp_510, while_asn_25_itm_1);
  assign and_347_nl = if_axi_wr_aw_PopNB_mioi_bawt & (~ mux_tmp_611);
  assign mux_612_nl = MUX_s_1_2_2(and_347_nl, and_tmp_71, if_axi_wr_aw_PopNB_mioi_ivld_mxwt);
  assign mux_613_nl = MUX_s_1_2_2(mux_612_nl, (~ mux_tmp_611), while_asn_30_itm_1);
  assign mux_tmp_614 = MUX_s_1_2_2(mux_613_nl, and_tmp_72, write_arb_req_sva);
  assign or_tmp_514 = or_tmp_349 | (~ mux_610_itm);
  assign and_tmp_78 = or_dcpl_2 & mux_tmp_614;
  assign nand_tmp_102 = ~(or_dcpl_3 & (~ mux_tmp_611));
  assign nand_tmp_103 = ~(regIn_PopNB_mioi_bawt & (~ nand_tmp_102));
  assign or_693_nl = if_axi_wr_aw_PopNB_mioi_ivld_mxwt | (~ if_axi_wr_aw_PopNB_mioi_bawt)
      | mux_tmp_611;
  assign mux_tmp_622 = MUX_s_1_2_2(or_693_nl, mux_tmp_611, while_asn_30_itm_1);
  assign mux_630_nl = MUX_s_1_2_2(and_tmp_76, (~ or_tmp_509), arb_next_1_1_sva);
  assign nand_105_nl = ~(select_mask_2_1_sva_1 & mux_630_nl);
  assign nor_120_nl = ~(regIn_PopNB_mioi_ivld_mxwt | (~ and_tmp_75));
  assign mux_628_nl = MUX_s_1_2_2(nor_120_nl, and_tmp_72, while_asn_34_itm_1);
  assign or_592_nl = regIn_arb_req_sva | (~ mux_628_nl);
  assign mux_629_nl = MUX_s_1_2_2((~ and_tmp_76), or_592_nl, arb_next_1_2_sva);
  assign or_593_nl = select_mask_2_1_sva_1 | mux_629_nl;
  assign mux_631_nl = MUX_s_1_2_2(nand_105_nl, or_593_nl, select_mask_2_1_sva_0);
  assign or_590_nl = or_tmp_349 | mux_tmp_622;
  assign mux_623_nl = MUX_s_1_2_2(nand_tmp_103, or_590_nl, regIn_PopNB_mioi_ivld_mxwt);
  assign mux_624_nl = MUX_s_1_2_2(mux_623_nl, nand_tmp_102, while_asn_34_itm_1);
  assign or_588_nl = (~ or_dcpl_2) | write_arb_req_sva | mux_tmp_622;
  assign mux_625_nl = MUX_s_1_2_2(mux_624_nl, or_588_nl, regIn_arb_req_sva);
  assign mux_619_nl = MUX_s_1_2_2(nand_tmp_103, or_tmp_514, regIn_PopNB_mioi_ivld_mxwt);
  assign mux_620_nl = MUX_s_1_2_2(mux_619_nl, nand_tmp_102, while_asn_34_itm_1);
  assign mux_621_nl = MUX_s_1_2_2(mux_620_nl, or_tmp_509, regIn_arb_req_sva);
  assign mux_626_nl = MUX_s_1_2_2(mux_625_nl, mux_621_nl, arb_next_1_2_sva);
  assign nand_164_nl = ~(regIn_PopNB_mioi_bawt & mux_tmp_614);
  assign mux_615_nl = MUX_s_1_2_2(nand_164_nl, or_tmp_514, regIn_PopNB_mioi_ivld_mxwt);
  assign mux_616_nl = MUX_s_1_2_2(mux_615_nl, (~ mux_tmp_614), while_asn_34_itm_1);
  assign mux_617_nl = MUX_s_1_2_2(mux_616_nl, or_tmp_509, regIn_arb_req_sva);
  assign mux_618_nl = MUX_s_1_2_2((~ and_tmp_78), mux_617_nl, arb_next_1_2_sva);
  assign mux_627_nl = MUX_s_1_2_2(mux_626_nl, mux_618_nl, arb_next_1_1_sva);
  assign mux_tmp_633 = MUX_s_1_2_2(mux_631_nl, mux_627_nl, arb_needs_update_sva);
  assign mux_638_nl = MUX_s_1_2_2(and_tmp_75, (~ or_tmp_514), regIn_PopNB_mioi_ivld_mxwt);
  assign mux_639_nl = MUX_s_1_2_2(mux_638_nl, and_tmp_72, while_asn_34_itm_1);
  assign mux_640_nl = MUX_s_1_2_2((~ mux_639_nl), or_tmp_509, regIn_arb_req_sva);
  assign mux_tmp_642 = MUX_s_1_2_2((~ and_tmp_76), mux_640_nl, or_tmp_292);
  assign not_tmp_372 = or_dcpl_2 & (~ nand_tmp_102);
  assign mux_651_nl = MUX_s_1_2_2(not_tmp_372, and_tmp_78, arb_next_1_1_sva);
  assign mux_tmp_653 = MUX_s_1_2_2((~ mux_tmp_633), mux_651_nl, operator_3_false_3_operator_3_false_3_and_svs_1);
  assign not_tmp_373 = MUX_s_1_2_2((~ mux_tmp_653), mux_tmp_633, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_tmp_656 = MUX_s_1_2_2(mux_tmp_633, mux_tmp_642, operator_8_false_operator_8_false_nor_mdf_sva);
  assign or_tmp_529 = write_arb_req_sva | (~ nand_tmp_98);
  assign mux_679_nl = MUX_s_1_2_2(operator_3_false_3_operator_3_false_3_and_svs_1,
      and_352_cse, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_677_nl = MUX_s_1_2_2(operator_8_false_operator_8_false_nor_mdf_sva,
      nor_116_cse, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_680_nl = MUX_s_1_2_2(mux_679_nl, mux_677_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign and_dcpl_130 = ~((mux_680_nl & while_stage_v_1) | arb_needs_update_sva);
  assign mux_456_nl = MUX_s_1_2_2(and_tmp_32, (~ or_tmp_287), write_arb_req_sva);
  assign nor_123_nl = ~(write_arb_req_sva | read_arb_req_sva | and_dcpl_35);
  assign mux_457_nl = MUX_s_1_2_2(mux_456_nl, nor_123_nl, regIn_arb_req_sva);
  assign nand_89_nl = ~(arb_needs_update_sva & mux_457_nl);
  assign and_256_cse = MUX_s_1_2_2(nand_89_nl, mux_tmp_455, while_stage_v_1);
  assign or_tmp_576 = or_dcpl_25 & (~ while_stage_v_1) & (fsm_output[1]);
  assign if_axi_rd_r_Push_mioi_idat_67_4_mx0c1 = and_dcpl_26 & (while_if_4_acc_1_itm_16_1
      | while_if_4_aelse_acc_itm_16_1) & and_dcpl;
  assign or_527_nl = or_tmp_435 | and_dcpl_35;
  assign or_525_nl = nor_tmp_30 | (~ and_tmp_32);
  assign or_524_nl = or_tmp_439 | (~ and_tmp_32);
  assign mux_576_nl = MUX_s_1_2_2(or_525_nl, or_524_nl, arb_next_1_1_sva);
  assign mux_577_nl = MUX_s_1_2_2(or_527_nl, mux_576_nl, arb_needs_update_sva);
  assign mux_578_nl = MUX_s_1_2_2(mux_577_nl, mux_tmp_575, while_stage_v_1);
  assign operator_3_false_2_operator_3_false_2_and_svs_st_1_mx0c1 = ((~ mux_578_nl)
      & (fsm_output[1])) | ((~ mux_tmp_575) & while_stage_v_1);
  assign nor_131_nl = ~(or_dcpl_4 | (~ mux_tmp_364));
  assign mux_579_nl = MUX_s_1_2_2(mux_tmp_364, nor_131_nl, or_dcpl_3);
  assign mux_580_nl = MUX_s_1_2_2(mux_tmp_364, mux_579_nl, or_dcpl_2);
  assign mux_581_nl = MUX_s_1_2_2(mux_tmp_364, mux_580_nl, or_234_cse);
  assign mux_582_nl = MUX_s_1_2_2(mux_tmp_364, mux_581_nl, while_stage_v_1);
  assign while_stage_v_2_mx0c1 = mux_582_nl & while_stage_v_2;
  assign or_539_nl = (~ if_axi_wr_w_PopNB_mioi_bawt) | if_axi_wr_w_PopNB_mioi_ivld_mxwt
      | and_dcpl_35;
  assign mux_588_nl = MUX_s_1_2_2(and_dcpl_35, or_539_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_589_nl = MUX_s_1_2_2((~ mux_588_nl), or_dcpl_25, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1_mx0c1 =
      mux_589_nl & or_dcpl_4 & or_dcpl_3 & or_dcpl_2 & while_stage_v_1;
  assign while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1_mx0c1
      = and_dcpl_26 & or_tmp_385 & while_stage_v_1;
  assign nl_while_if_4_aelse_acc_nl = ({1'b1 , operator_33_true_return_15_0_sva})
      + conv_u2u_16_17({(~ axiRdAddr_15_3_sva_dfm_1_mx0) , (~ axiRdAddr_2_0_sva_dfm_1_mx1)})
      + 17'b00000000000000001;
  assign while_if_4_aelse_acc_nl = nl_while_if_4_aelse_acc_nl[16:0];
  assign while_if_4_aelse_acc_itm_16_1 = readslicef_17_1_16(while_if_4_aelse_acc_nl);
  assign nor_334_nl = ~((~ (regwr_addr_6_3_sva[3])) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2:0]!=3'b000));
  assign and_572_nl = while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_nor_6_itm_1 & (operator_17_true_return_1_3_0_sva_1[3]);
  assign mux_tmp = MUX_s_1_2_2(nor_334_nl, and_572_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nor_335_nl = ~((regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2:0]!=3'b100));
  assign and_573_nl = while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_nor_3_itm_1 & (operator_17_true_return_1_3_0_sva_1[2]);
  assign mux_tmp_683 = MUX_s_1_2_2(nor_335_nl, and_573_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign nor_336_nl = ~((~ operator_3_false_3_operator_3_false_3_and_svs_2) | (regwr_addr_6_3_sva!=4'b0010));
  assign and_574_nl = while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & (operator_17_true_return_1_3_0_sva_1[1]) & while_else_4_if_if_for_nor_1_itm_1;
  assign mux_tmp_686 = MUX_s_1_2_2(nor_336_nl, and_574_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_380_nl = nand_142_cse_1 & mux_tmp_686;
  assign and_379_nl = if_axi_rd_r_Push_mioi_bawt & mux_tmp_686;
  assign mux_tmp_687 = MUX_s_1_2_2(and_380_nl, and_379_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nor_tmp_73 = ((regwr_addr_6_3_sva!=4'b0010)) & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & (operator_17_true_return_1_3_0_sva_1[1]) & while_else_4_if_if_for_nor_1_itm_1;
  assign and_383_nl = nand_142_cse_1 & operator_3_false_2_operator_3_false_2_and_svs_2
      & nor_tmp_73;
  assign and_382_nl = if_axi_rd_r_Push_mioi_bawt & operator_3_false_2_operator_3_false_2_and_svs_2
      & nor_tmp_73;
  assign mux_tmp_688 = MUX_s_1_2_2(and_383_nl, and_382_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign and_dcpl_141 = run_wen & while_stage_v_2;
  assign nor_tmp_75 = while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & (operator_17_true_return_1_3_0_sva_1[0]) & while_else_4_if_if_for_nor_itm_1;
  assign nor_338_nl = ~((~ operator_3_false_3_operator_3_false_3_and_svs_2) | (regwr_addr_6_3_sva!=4'b0001));
  assign mux_tmp_696 = MUX_s_1_2_2(nor_338_nl, nor_tmp_75, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_390_nl = nand_142_cse_1 & mux_tmp_696;
  assign and_389_nl = if_axi_rd_r_Push_mioi_bawt & mux_tmp_696;
  assign mux_tmp_697 = MUX_s_1_2_2(and_390_nl, and_389_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nor_339_nl = ~((regwr_addr_6_3_sva[0]) | (~ nor_tmp_75));
  assign or_722_nl = (regwr_addr_6_3_sva[3:1]!=3'b000);
  assign mux_tmp_699 = MUX_s_1_2_2(nor_339_nl, nor_tmp_75, or_722_nl);
  assign and_392_nl = nand_142_cse_1 & operator_3_false_2_operator_3_false_2_and_svs_2
      & mux_tmp_699;
  assign and_391_nl = if_axi_rd_r_Push_mioi_bawt & operator_3_false_2_operator_3_false_2_and_svs_2
      & mux_tmp_699;
  assign mux_tmp_700 = MUX_s_1_2_2(and_392_nl, and_391_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign or_tmp_614 = and_515_cse | (~((~(and_512_cse | while_else_4_if_if_for_equal_tmp_3_1
      | while_else_4_if_if_for_equal_tmp_5_1 | while_else_4_if_if_for_equal_tmp_6_1
      | while_else_4_if_if_for_equal_tmp_7_1 | while_else_4_if_if_for_equal_tmp_9_1
      | while_else_4_if_if_for_equal_tmp_10_1 | while_else_4_if_if_for_equal_tmp_11_1
      | while_else_4_if_if_for_equal_tmp_12_1 | while_else_4_if_if_for_equal_tmp_13_1
      | while_else_4_if_if_for_while_else_4_if_if_for_and_13_itm_1 | while_else_4_if_if_for_while_else_4_if_if_for_and_14_itm_1
      | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)))
      & (~(and_517_cse | and_513_cse))));
  assign nand_tmp_110 = ~(operator_3_false_2_operator_3_false_2_and_svs_2 & (~ or_tmp_614));
  assign mux_tmp_708 = MUX_s_1_2_2((~ operator_3_false_3_operator_3_false_3_and_svs_2),
      or_tmp_614, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign or_730_nl = if_axi_wr_w_PopNB_mioi_bawt | (regwr_addr_6_3_sva!=4'b0000);
  assign mux_tmp_709 = MUX_s_1_2_2(mux_tmp_708, nand_tmp_110, or_730_nl);
  assign or_732_nl = (regwr_addr_6_3_sva!=4'b0000);
  assign mux_tmp_712 = MUX_s_1_2_2(mux_tmp_708, nand_tmp_110, or_732_nl);
  assign or_1052_nl = (~((regIn_PopNB_mioi_idat_mxwt[2:0]!=3'b000))) | mux_tmp_712;
  assign mux_718_nl = MUX_s_1_2_2(nand_tmp_110, or_1052_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_719_nl = MUX_s_1_2_2(mux_718_nl, mux_tmp_709, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_720_nl = MUX_s_1_2_2(mux_719_nl, nand_tmp_110, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_721_nl = MUX_s_1_2_2(mux_720_nl, mux_tmp_712, regIn_PopNB_mioi_idat_mxwt[3]);
  assign nand_180_nl = ~(((~ operator_3_false_3_operator_3_false_3_and_svs_st_1)
      | (regwr_addr_6_3_sva!=4'b0000)) & operator_3_false_2_operator_3_false_2_and_svs_2
      & (~ or_tmp_614));
  assign mux_715_nl = MUX_s_1_2_2(nand_180_nl, mux_tmp_709, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_716_nl = MUX_s_1_2_2(mux_715_nl, nand_tmp_110, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_722_nl = MUX_s_1_2_2(mux_721_nl, mux_716_nl, regIn_arb_req_sva);
  assign mux_723_nl = MUX_s_1_2_2(mux_tmp_712, mux_722_nl, or_dcpl_4);
  assign nor_160_nl = ~((~ or_dcpl_3) | (~ while_stage_v_1) | operator_3_false_1_operator_3_false_1_and_svs_1
      | operator_3_false_2_operator_3_false_2_and_svs_1 | (~ operator_3_false_3_operator_3_false_3_and_svs_1));
  assign mux_724_nl = MUX_s_1_2_2(mux_tmp_712, mux_723_nl, nor_160_nl);
  assign mux_725_itm = MUX_s_1_2_2(mux_tmp_712, mux_724_nl, or_dcpl_2);
  assign and_589_nl = nand_142_cse_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_9_1;
  assign and_590_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_9_1;
  assign mux_tmp_722 = MUX_s_1_2_2(and_589_nl, and_590_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nor_343_nl = ~(and_302_cse | (~ (regwr_addr_6_3_sva[3])) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2:0]!=3'b001));
  assign nor_344_nl = ~((~ if_axi_rd_r_Push_mioi_bawt) | (~ (regwr_addr_6_3_sva[3]))
      | (~ operator_3_false_3_operator_3_false_3_and_svs_2) | (regwr_addr_6_3_sva[2:0]!=3'b001));
  assign not_tmp_415 = MUX_s_1_2_2(nor_343_nl, nor_344_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_724 = MUX_s_1_2_2(not_tmp_415, mux_tmp_722, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign or_746_cse = (~ operator_3_false_2_operator_3_false_2_and_svs_1) | operator_3_false_1_operator_3_false_1_and_svs_st_1
      | operator_3_false_2_operator_3_false_2_and_svs_st_1;
  assign and_592_nl = or_746_cse & not_tmp_415;
  assign mux_730_itm = MUX_s_1_2_2(and_592_nl, mux_tmp_722, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_594_nl = nand_142_cse_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_10_1;
  assign and_595_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_10_1;
  assign mux_tmp_730 = MUX_s_1_2_2(and_594_nl, and_595_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nor_345_nl = ~(and_302_cse | (~ (regwr_addr_6_3_sva[3])) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2:0]!=3'b010));
  assign nor_346_nl = ~((~ if_axi_rd_r_Push_mioi_bawt) | (~ (regwr_addr_6_3_sva[3]))
      | (~ operator_3_false_3_operator_3_false_3_and_svs_2) | (regwr_addr_6_3_sva[2:0]!=3'b010));
  assign not_tmp_422 = MUX_s_1_2_2(nor_345_nl, nor_346_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_732 = MUX_s_1_2_2(not_tmp_422, mux_tmp_730, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_597_nl = or_746_cse & not_tmp_422;
  assign mux_738_itm = MUX_s_1_2_2(and_597_nl, mux_tmp_730, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_599_nl = nand_142_cse_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_6_1;
  assign and_600_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_6_1;
  assign mux_tmp_738 = MUX_s_1_2_2(and_599_nl, and_600_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nor_347_nl = ~(and_302_cse | (regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2:0]!=3'b110));
  assign nor_348_nl = ~((~ if_axi_rd_r_Push_mioi_bawt) | (regwr_addr_6_3_sva[3])
      | (~ operator_3_false_3_operator_3_false_3_and_svs_2) | (regwr_addr_6_3_sva[2:0]!=3'b110));
  assign not_tmp_429 = MUX_s_1_2_2(nor_347_nl, nor_348_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_740 = MUX_s_1_2_2(not_tmp_429, mux_tmp_738, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_602_nl = or_746_cse & not_tmp_429;
  assign mux_746_itm = MUX_s_1_2_2(and_602_nl, mux_tmp_738, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_604_nl = nand_142_cse_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_11_1;
  assign and_605_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_11_1;
  assign mux_tmp_746 = MUX_s_1_2_2(and_604_nl, and_605_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign not_tmp_436 = ~((regwr_addr_6_3_sva[1:0]==2'b11));
  assign nor_349_nl = ~(and_302_cse | (~ (regwr_addr_6_3_sva[3])) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2]) | not_tmp_436);
  assign nor_350_nl = ~((~(if_axi_rd_r_Push_mioi_bawt & (regwr_addr_6_3_sva[3]) &
      operator_3_false_3_operator_3_false_3_and_svs_2 & (~ (regwr_addr_6_3_sva[2]))))
      | not_tmp_436);
  assign not_tmp_437 = MUX_s_1_2_2(nor_349_nl, nor_350_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_748 = MUX_s_1_2_2(not_tmp_437, mux_tmp_746, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_608_nl = or_746_cse & not_tmp_437;
  assign mux_754_itm = MUX_s_1_2_2(and_608_nl, mux_tmp_746, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_610_nl = nand_142_cse_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_3_1;
  assign and_611_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_3_1;
  assign mux_tmp_754 = MUX_s_1_2_2(and_610_nl, and_611_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nor_351_nl = ~(and_302_cse | (regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2]) | not_tmp_436);
  assign nor_352_nl = ~((~ if_axi_rd_r_Push_mioi_bawt) | (regwr_addr_6_3_sva[3])
      | (~ operator_3_false_3_operator_3_false_3_and_svs_2) | (regwr_addr_6_3_sva[2])
      | not_tmp_436);
  assign not_tmp_445 = MUX_s_1_2_2(nor_351_nl, nor_352_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_756 = MUX_s_1_2_2(not_tmp_445, mux_tmp_754, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_614_nl = or_746_cse & not_tmp_445;
  assign mux_762_itm = MUX_s_1_2_2(and_614_nl, mux_tmp_754, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_616_nl = nand_142_cse_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_7_1;
  assign and_617_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_7_1;
  assign mux_tmp_762 = MUX_s_1_2_2(and_616_nl, and_617_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign not_tmp_452 = ~(operator_3_false_3_operator_3_false_3_and_svs_2 & (regwr_addr_6_3_sva[2:0]==3'b111));
  assign nor_353_nl = ~(and_302_cse | (regwr_addr_6_3_sva[3]) | not_tmp_452);
  assign nor_354_nl = ~((~ if_axi_rd_r_Push_mioi_bawt) | (regwr_addr_6_3_sva[3])
      | not_tmp_452);
  assign not_tmp_453 = MUX_s_1_2_2(nor_353_nl, nor_354_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_764 = MUX_s_1_2_2(not_tmp_453, mux_tmp_762, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_620_nl = or_746_cse & not_tmp_453;
  assign mux_770_itm = MUX_s_1_2_2(and_620_nl, mux_tmp_762, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_622_nl = nand_142_cse_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_12_1;
  assign and_623_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_12_1;
  assign mux_tmp_770 = MUX_s_1_2_2(and_622_nl, and_623_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nor_355_nl = ~(and_302_cse | (~ (regwr_addr_6_3_sva[3])) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2:0]!=3'b100));
  assign nor_356_nl = ~((~ if_axi_rd_r_Push_mioi_bawt) | (~ (regwr_addr_6_3_sva[3]))
      | (~ operator_3_false_3_operator_3_false_3_and_svs_2) | (regwr_addr_6_3_sva[2:0]!=3'b100));
  assign not_tmp_460 = MUX_s_1_2_2(nor_355_nl, nor_356_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_772 = MUX_s_1_2_2(not_tmp_460, mux_tmp_770, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_625_nl = or_746_cse & not_tmp_460;
  assign mux_778_itm = MUX_s_1_2_2(and_625_nl, mux_tmp_770, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_627_nl = nand_142_cse_1 & while_else_4_if_if_for_equal_tmp_13_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign and_628_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_if_for_equal_tmp_13_1
      & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1;
  assign mux_tmp_778 = MUX_s_1_2_2(and_627_nl, and_628_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign and_630_nl = nand_142_cse_1 & (regwr_addr_6_3_sva[3]) & operator_3_false_3_operator_3_false_3_and_svs_2
      & (regwr_addr_6_3_sva[2:0]==3'b101);
  assign and_631_nl = if_axi_rd_r_Push_mioi_bawt & (regwr_addr_6_3_sva[3]) & operator_3_false_3_operator_3_false_3_and_svs_2
      & (regwr_addr_6_3_sva[2:0]==3'b101);
  assign not_tmp_468 = MUX_s_1_2_2(and_630_nl, and_631_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_780 = MUX_s_1_2_2(not_tmp_468, mux_tmp_778, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_632_nl = or_746_cse & not_tmp_468;
  assign mux_786_itm = MUX_s_1_2_2(and_632_nl, mux_tmp_778, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_634_nl = nand_142_cse_1 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_5_1;
  assign and_635_nl = if_axi_rd_r_Push_mioi_bawt & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_5_1;
  assign mux_tmp_786 = MUX_s_1_2_2(and_634_nl, and_635_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nor_357_nl = ~(and_302_cse | (regwr_addr_6_3_sva[3]) | (~ operator_3_false_3_operator_3_false_3_and_svs_2)
      | (regwr_addr_6_3_sva[2:0]!=3'b101));
  assign nor_358_nl = ~((~ if_axi_rd_r_Push_mioi_bawt) | (regwr_addr_6_3_sva[3])
      | (~ operator_3_false_3_operator_3_false_3_and_svs_2) | (regwr_addr_6_3_sva[2:0]!=3'b101));
  assign not_tmp_476 = MUX_s_1_2_2(nor_357_nl, nor_358_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_tmp_788 = MUX_s_1_2_2(not_tmp_476, mux_tmp_786, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_637_nl = or_746_cse & not_tmp_476;
  assign mux_794_itm = MUX_s_1_2_2(and_637_nl, mux_tmp_786, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign or_tmp_728 = while_asn_25_itm_1 | (~ if_axi_rd_ar_PopNB_mioi_bawt);
  assign or_841_cse = (~ if_axi_rd_ar_PopNB_mioi_ivld_mxwt) | read_arb_req_sva;
  assign and_638_nl = ((if_axi_rd_ar_PopNB_mioi_idat_mxwt[27:20]!=8'b00000000)) &
      operator_3_false_1_operator_3_false_1_and_svs_1;
  assign mux_799_nl = MUX_s_1_2_2((~ or_tmp_728), or_dcpl_4, and_638_nl);
  assign and_436_nl = ((axiRdLen_sva!=8'b00000000)) & operator_3_false_1_operator_3_false_1_and_svs_1
      & or_dcpl_4;
  assign mux_tmp_795 = MUX_s_1_2_2(mux_799_nl, and_436_nl, or_841_cse);
  assign not_tmp_484 = ~(while_stage_v_2 | (~ mux_tmp_795));
  assign mux_802_nl = MUX_s_1_2_2(or_tmp_728, (~ or_dcpl_4), operator_3_false_1_operator_3_false_1_and_svs_1);
  assign mux_803_nl = MUX_s_1_2_2(mux_802_nl, or_tmp_728, operator_8_false_operator_8_false_nor_mdf_sva);
  assign or_849_nl = operator_8_false_operator_8_false_nor_mdf_sva | (~(operator_3_false_1_operator_3_false_1_and_svs_1
      & or_dcpl_4));
  assign mux_804_nl = MUX_s_1_2_2(mux_803_nl, or_849_nl, or_841_cse);
  assign nand_tmp_124 = (~((~ operator_3_false_2_operator_3_false_2_and_svs_st_1)
      | if_axi_wr_w_PopNB_mioi_bawt)) | mux_804_nl;
  assign and_dcpl_196 = if_axi_wr_w_PopNB_mioi_ivld_mxwt & operator_3_false_2_operator_3_false_2_and_svs_st_1;
  assign nor_tmp_125 = (operator_17_true_return_1_3_0_sva_1[3]) & while_else_4_if_if_for_nor_6_itm_1
      & (while_else_4_if_if_regAddr_acc_itm_6_3[3]);
  assign nor_367_nl = ~(and_512_cse | while_else_4_if_if_for_equal_tmp_12_1 | and_517_cse
      | while_else_4_if_if_for_equal_tmp_10_1 | (while_else_4_if_if_regAddr_acc_itm_6_3[3]));
  assign mux_828_nl = MUX_s_1_2_2(nor_367_nl, (while_else_4_if_if_regAddr_acc_itm_6_3[3]),
      and_515_cse);
  assign or_880_nl = while_else_4_if_if_for_while_else_4_if_if_for_and_13_itm_1 |
      while_else_4_if_if_for_while_else_4_if_if_for_and_14_itm_1 | while_else_4_if_if_for_equal_tmp_13_1
      | while_else_4_if_if_for_equal_tmp_11_1 | while_else_4_if_if_for_equal_tmp_9_1
      | while_else_4_if_if_for_equal_tmp_7_1 | while_else_4_if_if_for_equal_tmp_6_1
      | while_else_4_if_if_for_equal_tmp_5_1 | while_else_4_if_if_for_equal_tmp_3_1;
  assign mux_829_nl = MUX_s_1_2_2(mux_828_nl, nor_tmp_125, or_880_nl);
  assign and_646_nl = while_else_4_if_if_for_equal_tmp_9_1 & (while_else_4_if_if_regAddr_acc_itm_6_3[3]);
  assign mux_830_nl = MUX_s_1_2_2(mux_829_nl, and_646_nl, while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign or_879_nl = while_else_4_if_if_for_equal_tmp_9_1 | (~ (while_else_4_if_if_regAddr_acc_itm_6_3[3]));
  assign mux_827_nl = MUX_s_1_2_2(nor_tmp_125, or_879_nl, while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign mux_831_nl = MUX_s_1_2_2(mux_830_nl, mux_827_nl, and_513_cse);
  assign and_648_nl = while_else_4_if_if_for_equal_tmp_12_1 & (while_else_4_if_if_regAddr_acc_itm_6_3[3]);
  assign or_878_nl = while_else_4_if_if_for_equal_tmp_12_1 | (~ (while_else_4_if_if_regAddr_acc_itm_6_3[3]));
  assign mux_825_nl = MUX_s_1_2_2(and_648_nl, or_878_nl, and_512_cse);
  assign nor_368_nl = ~((~ while_else_4_if_if_for_equal_tmp_5_1) | (while_else_4_if_if_regAddr_acc_itm_6_3[3]));
  assign mux_824_nl = MUX_s_1_2_2(nor_368_nl, or_1037_cse, while_else_4_if_if_for_equal_tmp_13_1);
  assign mux_826_nl = MUX_s_1_2_2(mux_825_nl, mux_824_nl, while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign mux_832_nl = MUX_s_1_2_2(mux_831_nl, mux_826_nl, while_else_4_if_if_regAddr_acc_itm_6_3[2]);
  assign nand_277_nl = ~(while_else_4_if_if_for_equal_tmp_10_1 & (while_else_4_if_if_regAddr_acc_itm_6_3[3]));
  assign nor_370_nl = ~(while_else_4_if_if_for_equal_tmp_10_1 | (~ (while_else_4_if_if_regAddr_acc_itm_6_3[3])));
  assign mux_821_nl = MUX_s_1_2_2(nand_277_nl, nor_370_nl, and_517_cse);
  assign or_1060_nl = (~ while_else_4_if_if_for_equal_tmp_3_1) | (while_else_4_if_if_regAddr_acc_itm_6_3[3]);
  assign nor_371_nl = ~(while_else_4_if_if_for_equal_tmp_3_1 | (while_else_4_if_if_regAddr_acc_itm_6_3[3]));
  assign mux_820_nl = MUX_s_1_2_2(or_1060_nl, nor_371_nl, while_else_4_if_if_for_equal_tmp_11_1);
  assign mux_822_nl = MUX_s_1_2_2(mux_821_nl, mux_820_nl, while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign or_872_nl = (~ while_else_4_if_if_for_equal_tmp_6_1) | (while_else_4_if_if_regAddr_acc_itm_6_3[3]);
  assign or_871_nl = (~ while_else_4_if_if_for_equal_tmp_7_1) | (while_else_4_if_if_regAddr_acc_itm_6_3[3]);
  assign mux_819_nl = MUX_s_1_2_2(or_872_nl, or_871_nl, while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign mux_823_nl = MUX_s_1_2_2(mux_822_nl, mux_819_nl, while_else_4_if_if_regAddr_acc_itm_6_3[2]);
  assign mux_833_cse = MUX_s_1_2_2((~ mux_832_nl), mux_823_nl, while_else_4_if_if_regAddr_acc_itm_6_3[1]);
  assign or_tmp_762 = operator_3_false_1_operator_3_false_1_and_svs_2 | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ operator_3_false_2_operator_3_false_2_and_svs_2) | (~ while_else_4_if_if_while_else_4_if_if_nand_tmp_1)
      | (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[2]) | mux_833_cse;
  assign or_tmp_778 = operator_3_false_1_operator_3_false_1_and_svs_2 | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ operator_3_false_2_operator_3_false_2_and_svs_2) | (~ while_else_4_if_if_while_else_4_if_if_nand_tmp_1)
      | (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[1]) | mux_833_cse;
  assign or_tmp_794 = operator_3_false_1_operator_3_false_1_and_svs_2 | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ operator_3_false_2_operator_3_false_2_and_svs_2) | (~ while_else_4_if_if_while_else_4_if_if_nand_tmp_1)
      | (if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70[0]) | mux_833_cse;
  assign nor_tmp_150 = while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  assign not_tmp_533 = ~((while_else_4_if_if_regAddr_acc_itm_6_3[3]) | (~ nor_tmp_150));
  assign nor_tmp_158 = (operator_17_true_return_1_3_0_sva_1[3]) & while_else_4_if_if_for_nor_6_itm_1
      & (while_else_4_if_if_regAddr_acc_itm_6_3[3]) & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_while_else_4_if_if_nand_tmp_1;
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_b_Push_mioi_idat_3_0 <= 4'b0000;
    end
    else if ( if_axi_wr_bwrite_and_cse & ((and_dcpl_26 & write_arb_req_sva & if_axi_wr_w_PopNB_mioi_ivld_mxwt
        & and_dcpl_20 & and_dcpl_19) | and_44_rgt) ) begin
      if_axi_wr_b_Push_mioi_idat_3_0 <= MUX_v_4_2_2(axi_wr_req_addr_id_sva, (if_axi_wr_aw_PopNB_mioi_idat_mxwt[3:0]),
          and_44_rgt);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_b_Push_mioi_idat_5 <= 1'b0;
    end
    else if ( run_wen & (~(and_dcpl_35 | and_dcpl_34 | and_dcpl_33 | and_dcpl_32
        | (~(if_axi_wr_w_PopNB_mioi_ivld_mxwt & (if_axi_wr_w_PopNB_mioi_idat_mxwt[64])))
        | or_dcpl_28)) ) begin
      if_axi_wr_b_Push_mioi_idat_5 <= (z_out[16]) | (readslicef_17_1_16(while_else_4_if_if_acc_1_nl));
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_rd_r_Push_mioi_idat_3_0 <= 4'b0000;
    end
    else if ( if_axi_wr_bwrite_and_cse & ((and_dcpl_26 & read_arb_req_sva & operator_3_false_1_operator_3_false_1_and_svs_st_1
        & while_stage_v_1) | and_54_rgt) ) begin
      if_axi_rd_r_Push_mioi_idat_3_0 <= MUX_v_4_2_2(axi_rd_req_id_sva, (if_axi_rd_ar_PopNB_mioi_idat_mxwt[3:0]),
          and_54_rgt);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_rd_r_Push_mioi_idat_67_4 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((and_dcpl_26 & nor_124_cse & and_dcpl) | if_axi_rd_r_Push_mioi_idat_67_4_mx0c1)
        ) begin
      if_axi_rd_r_Push_mioi_idat_67_4 <= MUX_v_64_2_2(axi_rd_resp_data_sva_2, axi_rd_resp_data_sva,
          if_axi_rd_r_Push_mioi_idat_67_4_mx0c1);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_rd_r_Push_mioi_idat_69 <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_39) ) begin
      if_axi_rd_r_Push_mioi_idat_69 <= ~ nor_124_cse;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_rd_r_Push_mioi_idat_70 <= 1'b0;
    end
    else if ( if_axi_wr_bwrite_and_cse & (~ or_dcpl_39) ) begin
      if_axi_rd_r_Push_mioi_idat_70 <= operator_8_false_operator_8_false_nor_mdf_sva_mx1w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_b_Push_mioi_iswt0 <= 1'b0;
      if_axi_wr_w_PopNB_mioi_iswt0 <= 1'b0;
      if_axi_rd_r_Push_mioi_iswt0 <= 1'b0;
      regIn_PopNB_mioi_iswt0 <= 1'b0;
      if_axi_wr_aw_PopNB_mioi_iswt0 <= 1'b0;
      if_axi_rd_ar_PopNB_mioi_iswt0 <= 1'b0;
    end
    else if ( run_wen ) begin
      if_axi_wr_b_Push_mioi_iswt0 <= and_dcpl_26 & if_axi_wr_w_PopNB_mioi_ivld_mxwt
          & (if_axi_wr_w_PopNB_mioi_idat_mxwt[64]) & if_axi_wr_w_PopNB_mioi_bawt
          & and_dcpl_19;
      if_axi_wr_w_PopNB_mioi_iswt0 <= (~ mux_396_nl) & (fsm_output[1]);
      if_axi_rd_r_Push_mioi_iswt0 <= and_dcpl_26 & and_dcpl;
      regIn_PopNB_mioi_iswt0 <= (~ mux_403_nl) & (fsm_output[1]);
      if_axi_wr_aw_PopNB_mioi_iswt0 <= mux_411_nl & (fsm_output[1]);
      if_axi_rd_ar_PopNB_mioi_iswt0 <= (~ mux_417_nl) & (fsm_output[1]);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regOut_13 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_12 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_11 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_10 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_9 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_7 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_6 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_5 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      regOut_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( regOut_13_and_cse ) begin
      regOut_13 <= reg_13_sva_dfm_4_mx0w0;
      regOut_12 <= reg_12_sva_dfm_4_mx0w0;
      regOut_11 <= reg_11_sva_dfm_4_mx0w0;
      regOut_10 <= reg_10_sva_dfm_4_mx0w0;
      regOut_9 <= reg_9_sva_dfm_4_mx0w0;
      regOut_7 <= reg_7_sva_dfm_4_mx0w0;
      regOut_6 <= reg_6_sva_dfm_4_mx0w0;
      regOut_5 <= reg_5_sva_dfm_4_mx0w0;
      regOut_3 <= reg_3_sva_dfm_4_mx0w0;
      regOut_2 <= reg_2_sva_dfm_4_mx0w0;
      regOut_1 <= reg_1_sva_dfm_4_mx0w0;
      regOut_0 <= reg_0_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_regOut_8_cse <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_687_nl & (~ operator_3_false_1_operator_3_false_1_and_svs_2) &
        while_stage_v_2 & run_wen ) begin
      reg_regOut_8_cse <= reg_8_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_regOut_4_cse <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_690_nl & (~ operator_3_false_1_operator_3_false_1_and_svs_2) &
        while_stage_v_2 & run_wen ) begin
      reg_regOut_4_cse <= reg_4_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_2_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_700_nl & (~ (fsm_output[0])) & run_wen & (~ operator_3_false_1_operator_3_false_1_and_svs_2)
        & while_stage_v_2 ) begin
      reg_2_sva <= reg_2_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_1_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_712_nl & nor_303_cse & and_dcpl_141 ) begin
      reg_1_sva <= reg_1_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_0_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_726_nl & nor_303_cse & and_dcpl_141 ) begin
      reg_0_sva <= reg_0_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_9_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_734_nl & (~ operator_3_false_1_operator_3_false_1_and_svs_2) &
        while_stage_v_2 & (~ (fsm_output[0])) & run_wen ) begin
      reg_9_sva <= reg_9_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_10_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_742_nl & nor_303_cse & and_dcpl_141 ) begin
      reg_10_sva <= reg_10_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_6_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_750_nl & nor_303_cse & and_dcpl_141 ) begin
      reg_6_sva <= reg_6_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_11_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_758_nl & (~ operator_3_false_1_operator_3_false_1_and_svs_2) &
        while_stage_v_2 & (~ (fsm_output[0])) & run_wen ) begin
      reg_11_sva <= reg_11_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_3_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_766_nl & (~ operator_3_false_1_operator_3_false_1_and_svs_2) &
        while_stage_v_2 & (~ (fsm_output[0])) & run_wen ) begin
      reg_3_sva <= reg_3_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_7_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_774_nl & (~ operator_3_false_1_operator_3_false_1_and_svs_2) &
        while_stage_v_2 & (~ (fsm_output[0])) & run_wen ) begin
      reg_7_sva <= reg_7_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_12_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_782_nl & nor_303_cse & and_dcpl_141 ) begin
      reg_12_sva <= reg_12_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_13_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_790_nl & (~ operator_3_false_1_operator_3_false_1_and_svs_2) &
        while_stage_v_2 & (~ (fsm_output[0])) & run_wen ) begin
      reg_13_sva <= reg_13_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      reg_5_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( mux_798_nl & (~ operator_3_false_1_operator_3_false_1_and_svs_2) &
        while_stage_v_2 & (~ (fsm_output[0])) & run_wen ) begin
      reg_5_sva <= reg_5_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm
          <= 1'b0;
    end
    else if ( run_wen & (~(and_256_cse | ((mux_tmp_455 | (~ while_stage_v_1)) & (fsm_output[0]))))
        ) begin
      nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm
          <= nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_0_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm
          <= 1'b0;
      arb_pick_if_1_and_tmp_2 <= 1'b0;
      arb_pick_if_1_and_stg_1_0 <= 1'b0;
      arb_pick_priority_4_sva <= 1'b0;
      operator_5_false_operator_5_false_operator_5_false_or_svs <= 1'b0;
    end
    else if ( nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_and_1_cse
        ) begin
      nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm
          <= nvhls_leading_ones_5U_Arbiter_3U_Roundrobin_UnrolledMask_nvhls_nvhls_t_3U_nvuint_t_idx_1_lpi_1_dfm_mx0w0;
      arb_pick_if_1_and_tmp_2 <= arb_pick_if_1_and_tmp_2_mx0w0;
      arb_pick_if_1_and_stg_1_0 <= arb_pick_if_1_and_stg_1_0_mx0w0;
      arb_pick_priority_4_sva <= arb_pick_priority_4_sva_mx0w0;
      operator_5_false_operator_5_false_operator_5_false_or_svs <= operator_5_false_operator_5_false_operator_5_false_or_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regIn_arb_req_sva <= 1'b0;
      read_arb_req_sva <= 1'b0;
      write_arb_req_sva <= 1'b0;
    end
    else if ( regIn_arb_req_and_cse ) begin
      regIn_arb_req_sva <= MUX_s_1_2_2(while_while_or_2_tmp, while_else_4_mux_20_nl,
          and_dcpl_81);
      read_arb_req_sva <= MUX_s_1_2_2(while_if_4_while_if_4_and_1_mx0w0, while_while_or_tmp,
          and_dcpl_81);
      write_arb_req_sva <= MUX_s_1_2_2(while_while_or_1_tmp, while_else_4_mux_22_nl,
          and_dcpl_81);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      arb_next_1_2_sva <= 1'b1;
      arb_next_1_1_sva <= 1'b1;
    end
    else if ( arb_next_and_cse ) begin
      arb_next_1_2_sva <= arb_pick_if_1_not_15;
      arb_next_1_1_sva <= nvhls_set_slc_Arbiter_3U_Roundrobin_Mask_nvhls_nvhls_t_2U_nvuint_t_X_temp_2_1_sva_1_1
          | arb_pick_if_1_not_15;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      select_mask_0_sva <= 1'b0;
      select_mask_2_1_sva_1 <= 1'b0;
      select_mask_2_1_sva_0 <= 1'b0;
    end
    else if ( select_mask_and_cse ) begin
      select_mask_0_sva <= arb_pick_return_0_lpi_1_dfm_2;
      select_mask_2_1_sva_1 <= arb_pick_return_2_1_lpi_1_dfm_1_1_1;
      select_mask_2_1_sva_0 <= arb_pick_return_2_1_lpi_1_dfm_1_0_1;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      arb_needs_update_sva <= 1'b1;
      while_stage_v_1 <= 1'b0;
      operator_3_false_1_operator_3_false_1_and_svs_st_1 <= 1'b0;
    end
    else if ( arb_needs_update_and_cse ) begin
      arb_needs_update_sva <= (~(arb_pick_return_2_1_lpi_1_dfm_1_1_1 | arb_pick_return_2_1_lpi_1_dfm_1_0_1
          | arb_pick_return_0_lpi_1_dfm_2)) & while_if_4_mux1h_3_nl;
      while_stage_v_1 <= 1'b1;
      operator_3_false_1_operator_3_false_1_and_svs_st_1 <= operator_3_false_1_operator_3_false_1_and_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      axiRdAddr_2_0_sva_dfm_1 <= 3'b000;
    end
    else if ( run_wen & (~(while_asn_25_itm_1 | (~(if_axi_rd_ar_PopNB_mioi_ivld_mxwt
        & if_axi_rd_ar_PopNB_mioi_bawt & or_dcpl_25)) | or_dcpl_36 | and_dcpl_83
        | read_arb_req_sva | (~ while_stage_v_1))) ) begin
      axiRdAddr_2_0_sva_dfm_1 <= if_axi_rd_ar_PopNB_mioi_idat_mxwt[6:4];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      axiRdAddr_15_3_sva <= 13'b0000000000000;
      axiRdLen_sva <= 8'b00000000;
    end
    else if ( and_440_cse ) begin
      axiRdAddr_15_3_sva <= MUX_v_13_2_2(z_out_1, axiRdAddr_15_3_sva_dfm_1_mx0, and_dcpl_91);
      axiRdLen_sva <= MUX_v_8_2_2(while_if_4_else_2_acc_nl, axiRdLen_sva_dfm_1_mx0,
          and_dcpl_91);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      axiWrAddr_2_0_sva_dfm_1 <= 3'b000;
    end
    else if ( if_axi_wr_bwrite_and_cse & (~(or_tmp_282 | (~(if_axi_wr_aw_PopNB_mioi_bawt
        & or_dcpl_25)) | and_dcpl_34 | and_dcpl_32 | and_dcpl_83 | write_arb_req_sva
        | (~ while_stage_v_1))) ) begin
      axiWrAddr_2_0_sva_dfm_1 <= if_axi_wr_aw_PopNB_mioi_idat_mxwt[6:4];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      axiWrAddr_15_3_sva <= 13'b0000000000000;
    end
    else if ( run_wen & ((mux_501_nl & or_dcpl_4 & or_dcpl_3 & or_dcpl_2 & operator_3_false_2_operator_3_false_2_and_svs_1
        & (~ operator_3_false_1_operator_3_false_1_and_svs_1) & while_stage_v_1)
        | while_and_rgt) ) begin
      axiWrAddr_15_3_sva <= MUX_v_13_2_2(z_out_1, (if_axi_wr_aw_PopNB_mioi_idat_mxwt[19:7]),
          while_and_rgt);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_8_false_operator_8_false_nor_mdf_sva <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_35) ) begin
      operator_8_false_operator_8_false_nor_mdf_sva <= operator_8_false_operator_8_false_nor_mdf_sva_mx1w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      axi_rd_resp_data_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(mux_506_nl | and_dcpl_34 | or_dcpl_36 | (~(operator_3_false_1_operator_3_false_1_and_svs_1
        & while_stage_v_1)))) ) begin
      axi_rd_resp_data_sva <= axi_rd_resp_data_sva_2;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_33_true_return_15_0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (~ (fsm_output[1])) ) begin
      operator_33_true_return_15_0_sva <= z_out[15:0];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_3_false_2_operator_3_false_2_and_svs_st_1 <= 1'b0;
    end
    else if ( run_wen & ((mux_550_nl & (fsm_output[1])) | (mux_tmp_545 & while_stage_v_1)
        | operator_3_false_2_operator_3_false_2_and_svs_st_1_mx0c1) ) begin
      operator_3_false_2_operator_3_false_2_and_svs_st_1 <= MUX_s_1_2_2(operator_3_false_2_operator_3_false_2_and_svs_mx0w0,
          operator_3_false_2_operator_3_false_2_and_svs_st, operator_3_false_2_operator_3_false_2_and_svs_st_1_mx0c1);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_3_false_3_operator_3_false_3_and_svs_1 <= 1'b0;
      operator_3_false_2_operator_3_false_2_and_svs_1 <= 1'b0;
      operator_3_false_1_operator_3_false_1_and_svs_1 <= 1'b0;
    end
    else if ( operator_3_false_3_and_cse ) begin
      operator_3_false_3_operator_3_false_3_and_svs_1 <= operator_3_false_3_operator_3_false_3_and_svs_mx0w0;
      operator_3_false_2_operator_3_false_2_and_svs_1 <= operator_3_false_2_operator_3_false_2_and_svs_mx0w0;
      operator_3_false_1_operator_3_false_1_and_svs_1 <= operator_3_false_1_operator_3_false_1_and_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      axi_wr_req_addr_id_sva <= 4'b0000;
    end
    else if ( run_wen & (~ write_arb_req_sva) ) begin
      axi_wr_req_addr_id_sva <= if_axi_wr_aw_PopNB_mioi_idat_mxwt[3:0];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      axi_rd_req_id_sva <= 4'b0000;
    end
    else if ( run_wen & (~ read_arb_req_sva) ) begin
      axi_rd_req_id_sva <= if_axi_rd_ar_PopNB_mioi_idat_mxwt[3:0];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_asn_34_itm_1 <= 1'b0;
      while_asn_30_itm_1 <= 1'b0;
      while_asn_25_itm_1 <= 1'b0;
    end
    else if ( while_and_98_cse ) begin
      while_asn_34_itm_1 <= MUX1HOT_s_1_3_2(while_while_or_2_tmp, while_else_4_else_while_else_4_else_and_itm,
          regIn_arb_req_sva, {while_or_25_nl , while_and_103_cse , or_tmp_576});
      while_asn_30_itm_1 <= MUX1HOT_s_1_3_2(while_while_or_1_tmp, while_else_4_if_if_while_else_4_if_if_and_1_itm,
          write_arb_req_sva, {while_or_26_nl , while_and_108_nl , or_tmp_576});
      while_asn_25_itm_1 <= MUX1HOT_s_1_3_2(while_if_4_while_if_4_and_1_mx0w0, while_while_or_tmp,
          read_arb_req_sva, {and_dcpl_79 , and_dcpl_81 , or_tmp_576});
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_stage_v_2 <= 1'b0;
    end
    else if ( run_wen & ((and_dcpl_78 & while_stage_v_1) | while_stage_v_2_mx0c1)
        ) begin
      while_stage_v_2 <= ~ while_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1 <= 1'b0;
    end
    else if ( run_wen & ((and_dcpl_26 & if_axi_wr_w_PopNB_mioi_ivld_mxwt & if_axi_wr_w_PopNB_mioi_bawt
        & operator_3_false_2_operator_3_false_2_and_svs_st_1 & and_dcpl_55) | while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1_mx0c1)
        ) begin
      while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1 <= MUX_s_1_2_2((if_axi_wr_w_PopNB_mioi_idat_mxwt[64]),
          while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm, while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1_mx0c1);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_17_true_return_1_3_0_sva_1 <= 4'b0000;
      while_else_4_if_if_for_nor_6_itm_1 <= 1'b0;
      while_else_4_if_if_for_nor_3_itm_1 <= 1'b0;
      while_else_4_if_if_for_nor_1_itm_1 <= 1'b0;
      while_else_4_if_if_for_nor_itm_1 <= 1'b0;
    end
    else if ( while_else_4_if_if_regAddr_and_1_cse ) begin
      operator_17_true_return_1_3_0_sva_1 <= while_else_4_if_if_regAddr_acc_itm_6_3;
      while_else_4_if_if_for_nor_6_itm_1 <= ~((while_else_4_if_if_regAddr_acc_itm_6_3[2:0]!=3'b000));
      while_else_4_if_if_for_nor_3_itm_1 <= ~((while_else_4_if_if_regAddr_acc_itm_6_3[3])
          | (while_else_4_if_if_regAddr_acc_itm_6_3[1]) | (while_else_4_if_if_regAddr_acc_itm_6_3[0]));
      while_else_4_if_if_for_nor_1_itm_1 <= ~((while_else_4_if_if_regAddr_acc_itm_6_3[3])
          | (while_else_4_if_if_regAddr_acc_itm_6_3[2]) | (while_else_4_if_if_regAddr_acc_itm_6_3[0]));
      while_else_4_if_if_for_nor_itm_1 <= ~((while_else_4_if_if_regAddr_acc_itm_6_3[3:1]!=3'b000));
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~ mux_335_nl) & (~ and_dcpl_117) ) begin
      if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_63_0 <= if_axi_wr_w_PopNB_mioi_idat_mxwt[63:0];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_while_else_4_if_if_nand_tmp_1 <= 1'b0;
      if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70 <= 3'b000;
    end
    else if ( while_else_4_if_if_and_13_cse ) begin
      while_else_4_if_if_while_else_4_if_if_nand_tmp_1 <= ~((if_axi_wr_w_PopNB_mioi_idat_mxwt[72:65]==8'b11111111));
      if_axi_wr_w_PopNB_mio_mrgout_dat_sva_1_72_70 <= if_axi_wr_w_PopNB_mioi_idat_mxwt[72:70];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_if_1_for_8_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_63_56_itm_1
          <= 8'b00000000;
    end
    else if ( (~(mux_834_nl & while_stage_v_2)) & or_dcpl_3 & or_dcpl_2 & or_dcpl_4
        & if_axi_wr_w_PopNB_mioi_bawt & (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[72]))
        & run_wen & and_dcpl_196 & (~ operator_3_false_1_operator_3_false_1_and_svs_st_1)
        & operator_3_false_2_operator_3_false_2_and_svs_1 & (~ operator_3_false_1_operator_3_false_1_and_svs_1)
        & while_stage_v_1 ) begin
      while_else_4_if_if_if_1_for_8_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_63_56_itm_1
          <= while_else_4_if_if_if_1_old_data_sva_1[63:56];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_63_40 <= 24'b000000000000000000000000;
    end
    else if ( run_wen & (~ and_dcpl_117) ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_63_40 <= if_axi_wr_w_PopNB_mioi_idat_mxwt[63:40];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_if_1_for_7_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_55_48_itm_1
          <= 8'b00000000;
    end
    else if ( (~(mux_850_nl & while_stage_v_2)) & or_dcpl_3 & or_dcpl_2 & or_dcpl_4
        & if_axi_wr_w_PopNB_mioi_bawt & (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[71]))
        & run_wen & and_dcpl_196 & (~ operator_3_false_1_operator_3_false_1_and_svs_st_1)
        & operator_3_false_2_operator_3_false_2_and_svs_1 & (~ operator_3_false_1_operator_3_false_1_and_svs_1)
        & while_stage_v_1 ) begin
      while_else_4_if_if_if_1_for_7_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_55_48_itm_1
          <= while_else_4_if_if_if_1_old_data_sva_1[55:48];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_if_1_for_6_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_47_40_itm_1
          <= 8'b00000000;
    end
    else if ( (~(mux_866_nl & while_stage_v_2)) & or_dcpl_3 & or_dcpl_2 & or_dcpl_4
        & if_axi_wr_w_PopNB_mioi_bawt & (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[70]))
        & run_wen & and_dcpl_196 & (~ operator_3_false_1_operator_3_false_1_and_svs_st_1)
        & operator_3_false_2_operator_3_false_2_and_svs_1 & (~ operator_3_false_1_operator_3_false_1_and_svs_1)
        & while_stage_v_1 ) begin
      while_else_4_if_if_if_1_for_6_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_nvhls_get_slc_8U_nvhls_nvhls_t_64U_nvuint_t_slc_while_else_4_if_if_if_1_old_data_47_40_itm_1
          <= while_else_4_if_if_if_1_old_data_sva_1[47:40];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_39_32 <= 8'b00000000;
    end
    else if ( (~((~(or_927_cse & ((if_axi_wr_w_PopNB_mioi_idat_mxwt[69]) | (~ operator_3_false_2_operator_3_false_2_and_svs_2)
        | operator_3_false_1_operator_3_false_1_and_svs_2 | mux_884_cse))) & while_stage_v_2))
        & run_wen ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_39_32 <= MUX_v_8_2_2((if_axi_wr_w_PopNB_mioi_idat_mxwt[39:32]),
          (while_else_4_if_if_if_1_old_data_sva_1[39:32]), and_189_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_31_24 <= 8'b00000000;
    end
    else if ( (~((~(or_927_cse & ((if_axi_wr_w_PopNB_mioi_idat_mxwt[68]) | (~ operator_3_false_2_operator_3_false_2_and_svs_2)
        | operator_3_false_1_operator_3_false_1_and_svs_2 | mux_884_cse))) & while_stage_v_2))
        & run_wen ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_31_24 <= MUX_v_8_2_2((if_axi_wr_w_PopNB_mioi_idat_mxwt[31:24]),
          (while_else_4_if_if_if_1_old_data_sva_1[31:24]), and_191_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_23_16 <= 8'b00000000;
    end
    else if ( (~((~(or_927_cse & ((if_axi_wr_w_PopNB_mioi_idat_mxwt[67]) | (~ operator_3_false_2_operator_3_false_2_and_svs_2)
        | operator_3_false_1_operator_3_false_1_and_svs_2 | mux_884_cse))) & while_stage_v_2))
        & run_wen ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_23_16 <= MUX_v_8_2_2((if_axi_wr_w_PopNB_mioi_idat_mxwt[23:16]),
          (while_else_4_if_if_if_1_old_data_sva_1[23:16]), and_193_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_15_8 <= 8'b00000000;
    end
    else if ( (~((~(or_927_cse & ((if_axi_wr_w_PopNB_mioi_idat_mxwt[66]) | (~ operator_3_false_2_operator_3_false_2_and_svs_2)
        | operator_3_false_1_operator_3_false_1_and_svs_2 | mux_884_cse))) & while_stage_v_2))
        & run_wen ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_15_8 <= MUX_v_8_2_2((if_axi_wr_w_PopNB_mioi_idat_mxwt[15:8]),
          (while_else_4_if_if_if_1_old_data_sva_1[15:8]), and_195_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_7_0 <= 8'b00000000;
    end
    else if ( (~((~(or_927_cse & ((if_axi_wr_w_PopNB_mioi_idat_mxwt[65]) | (~ operator_3_false_2_operator_3_false_2_and_svs_2)
        | operator_3_false_1_operator_3_false_1_and_svs_2 | mux_884_cse))) & while_stage_v_2))
        & run_wen ) begin
      while_else_4_if_if_axiData_lpi_1_dfm_4_1_7_0 <= MUX_v_8_2_2((if_axi_wr_w_PopNB_mioi_idat_mxwt[7:0]),
          (while_else_4_if_if_if_1_old_data_sva_1[7:0]), and_197_nl);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
          <= 1'b0;
    end
    else if ( run_wen & (and_dcpl_58 | while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1_mx0c1)
        ) begin
      while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
          <= MUX_s_1_2_2(if_axi_wr_w_PopNB_mioi_ivld_mxwt, while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st,
          while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1_mx0c1);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_3_false_2_operator_3_false_2_and_svs_st_2 <= 1'b0;
      operator_3_false_1_operator_3_false_1_and_svs_st_2 <= 1'b0;
    end
    else if ( operator_3_false_2_and_2_cse ) begin
      operator_3_false_2_operator_3_false_2_and_svs_st_2 <= operator_3_false_2_operator_3_false_2_and_svs_st_1;
      operator_3_false_1_operator_3_false_1_and_svs_st_2 <= operator_3_false_1_operator_3_false_1_and_svs_st_1;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_3_false_1_operator_3_false_1_and_svs_2 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_13_1 <= 1'b0;
      while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
      operator_3_false_3_operator_3_false_3_and_svs_2 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_12_1 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_11_1 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_10_1 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_9_1 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_7_1 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_6_1 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_5_1 <= 1'b0;
      while_else_4_if_if_for_equal_tmp_3_1 <= 1'b0;
      operator_3_false_2_operator_3_false_2_and_svs_2 <= 1'b0;
      while_else_4_if_if_for_while_else_4_if_if_for_and_13_itm_1 <= 1'b0;
      while_else_4_if_if_for_while_else_4_if_if_for_and_14_itm_1 <= 1'b0;
    end
    else if ( operator_3_false_1_and_cse ) begin
      operator_3_false_1_operator_3_false_1_and_svs_2 <= operator_3_false_1_operator_3_false_1_and_svs_1;
      while_else_4_if_if_for_equal_tmp_13_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b1101);
      while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
          <= if_axi_wr_w_PopNB_mioi_ivld_mxwt;
      operator_3_false_3_operator_3_false_3_and_svs_2 <= operator_3_false_3_operator_3_false_3_and_svs_1;
      while_else_4_if_if_for_equal_tmp_12_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b1100);
      while_else_4_if_if_for_equal_tmp_11_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b1011);
      while_else_4_if_if_for_equal_tmp_10_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b1010);
      while_else_4_if_if_for_equal_tmp_9_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b1001);
      while_else_4_if_if_for_equal_tmp_7_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b0111);
      while_else_4_if_if_for_equal_tmp_6_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b0110);
      while_else_4_if_if_for_equal_tmp_5_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b0101);
      while_else_4_if_if_for_equal_tmp_3_1 <= (while_else_4_if_if_regAddr_acc_itm_6_3==4'b0011);
      operator_3_false_2_operator_3_false_2_and_svs_2 <= operator_3_false_2_operator_3_false_2_and_svs_1;
      while_else_4_if_if_for_while_else_4_if_if_for_and_13_itm_1 <= (operator_17_true_return_1_3_0_sva_mx1==4'b1110);
      while_else_4_if_if_for_while_else_4_if_if_for_and_14_itm_1 <= (operator_17_true_return_1_3_0_sva_mx1==4'b1111);
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      regwr_addr_6_3_sva <= 4'b0000;
      regwr_data_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( regwr_addr_and_cse ) begin
      regwr_addr_6_3_sva <= regIn_PopNB_mioi_idat_mxwt[3:0];
      regwr_data_sva <= regIn_PopNB_mioi_idat_mxwt[67:4];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_3_false_2_operator_3_false_2_and_svs_st <= 1'b0;
    end
    else if ( run_wen & (~ mux_675_nl) ) begin
      operator_3_false_2_operator_3_false_2_and_svs_st <= operator_3_false_2_operator_3_false_2_and_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_38 | or_dcpl_36 | (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt)
        | or_dcpl_28)) ) begin
      while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm <= if_axi_wr_w_PopNB_mioi_idat_mxwt[64];
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st
          <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_38 | or_dcpl_36 | or_dcpl_28)) ) begin
      while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st
          <= if_axi_wr_w_PopNB_mioi_ivld_mxwt;
    end
  end
  always @(posedge clk or negedge reset_bar) begin
    if ( ~ reset_bar ) begin
      operator_3_false_3_operator_3_false_3_and_svs_st_1 <= 1'b0;
    end
    else if ( run_wen & mux_676_nl ) begin
      operator_3_false_3_operator_3_false_3_and_svs_st_1 <= operator_3_false_3_operator_3_false_3_and_svs_mx0w0;
    end
  end
  assign nl_while_else_4_if_if_acc_1_nl = ({1'b1 , axiWrAddr_15_3_sva_dfm_1_mx0 ,
      axiWrAddr_2_0_sva_dfm_1_mx1}) + conv_u2u_16_17(~ baseAddr) + 17'b00000000000000001;
  assign while_else_4_if_if_acc_1_nl = nl_while_else_4_if_if_acc_1_nl[16:0];
  assign or_344_nl = or_tmp_280 | and_dcpl_35;
  assign or_342_nl = regIn_arb_req_sva | (~ write_arb_req_sva) | read_arb_req_sva
      | and_dcpl_35;
  assign or_340_nl = nor_tmp_30 | (~(write_arb_req_sva & or_dcpl_25));
  assign mux_394_nl = MUX_s_1_2_2(or_342_nl, or_340_nl, arb_next_1_1_sva);
  assign mux_395_nl = MUX_s_1_2_2(or_344_nl, mux_394_nl, arb_needs_update_sva);
  assign mux_391_nl = MUX_s_1_2_2(mux_682_itm, mux_tmp_378, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign or_337_nl = and_352_cse | mux_tmp_378;
  assign mux_389_nl = MUX_s_1_2_2(mux_682_itm, or_337_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nand_70_nl = ~(if_axi_wr_w_PopNB_mioi_bawt & (~ mux_389_nl));
  assign mux_392_nl = MUX_s_1_2_2(mux_391_nl, nand_70_nl, nor_tmp_28);
  assign nand_68_nl = ~(or_28_cse & (~ mux_tmp_378));
  assign nand_67_nl = ~(or_28_cse & (~ mux_tmp_381));
  assign mux_383_nl = MUX_s_1_2_2(nand_68_nl, nand_67_nl, operator_8_false_operator_8_false_nor_mdf_sva);
  assign mux_382_nl = MUX_s_1_2_2(mux_tmp_381, mux_tmp_378, or_310_cse);
  assign mux_384_nl = MUX_s_1_2_2(mux_383_nl, mux_382_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_393_nl = MUX_s_1_2_2(mux_392_nl, mux_384_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign mux_396_nl = MUX_s_1_2_2(mux_395_nl, mux_393_nl, while_stage_v_1);
  assign or_354_nl = regIn_arb_req_sva | (~ nand_tmp_71);
  assign nand_168_nl = ~(or_dcpl_2 & and_tmp_21);
  assign mux_399_nl = MUX_s_1_2_2(or_tmp_311, nand_168_nl, operator_3_false_3_operator_3_false_3_and_svs_1);
  assign or_347_nl = operator_3_false_1_operator_3_false_1_and_svs_1 | operator_3_false_2_operator_3_false_2_and_svs_1;
  assign mux_400_nl = MUX_s_1_2_2(mux_399_nl, or_tmp_311, or_347_nl);
  assign mux_401_nl = MUX_s_1_2_2(or_354_nl, mux_400_nl, while_stage_v_1);
  assign mux_402_nl = MUX_s_1_2_2(or_tmp_315, mux_401_nl, or_234_cse);
  assign mux_403_nl = MUX_s_1_2_2(or_tmp_315, mux_402_nl, or_dcpl_4);
  assign nor_125_nl = ~(write_arb_req_sva | and_dcpl_35);
  assign and_353_nl = operator_3_false_2_operator_3_false_2_and_svs_1 & (if_axi_wr_w_PopNB_mioi_idat_mxwt[64])
      & if_axi_wr_w_PopNB_mioi_ivld_mxwt;
  assign mux_406_nl = MUX_s_1_2_2((~ or_tmp_322), and_dcpl_26, and_353_nl);
  assign and_354_nl = if_axi_wr_w_PopNB_mioi_bawt & mux_406_nl;
  assign mux_409_nl = MUX_s_1_2_2((~ or_tmp_322), and_354_nl, nor_tmp_28);
  assign and_355_nl = or_234_cse & (~ or_tmp_322);
  assign mux_410_nl = MUX_s_1_2_2(mux_409_nl, and_355_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign mux_411_nl = MUX_s_1_2_2(nor_125_nl, mux_410_nl, while_stage_v_1);
  assign or_376_nl = read_arb_req_sva | (~ nand_tmp_71);
  assign mux_415_nl = MUX_s_1_2_2(not_tmp_258, nand_tmp_74, while_while_or_tmp);
  assign nand_75_nl = ~(if_axi_rd_ar_PopNB_mioi_bawt & (~ mux_415_nl));
  assign mux_414_nl = MUX_s_1_2_2(not_tmp_258, nand_tmp_74, read_arb_req_sva);
  assign mux_416_nl = MUX_s_1_2_2(nand_75_nl, mux_414_nl, while_asn_25_itm_1);
  assign mux_417_nl = MUX_s_1_2_2(or_376_nl, mux_416_nl, while_stage_v_1);
  assign and_501_nl = nand_198_cse & mux_tmp;
  assign mux_686_nl = MUX_s_1_2_2(and_501_nl, mux_tmp, if_axi_wr_b_Push_mioi_bawt);
  assign and_370_nl = if_axi_rd_r_Push_mioi_bawt & mux_tmp;
  assign mux_687_nl = MUX_s_1_2_2(mux_686_nl, and_370_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign and_503_nl = nand_198_cse & mux_tmp_683;
  assign mux_689_nl = MUX_s_1_2_2(and_503_nl, mux_tmp_683, if_axi_wr_b_Push_mioi_bawt);
  assign and_374_nl = if_axi_rd_r_Push_mioi_bawt & mux_tmp_683;
  assign mux_690_nl = MUX_s_1_2_2(mux_689_nl, and_374_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign and_384_nl = regIn_arb_req_sva & mux_tmp_688;
  assign mux_694_nl = MUX_s_1_2_2(mux_tmp_687, mux_tmp_688, regIn_arb_req_sva);
  assign or_710_nl = (regIn_PopNB_mioi_idat_mxwt[3:0]!=4'b0010);
  assign mux_695_nl = MUX_s_1_2_2(and_384_nl, mux_694_nl, or_710_nl);
  assign mux_696_nl = MUX_s_1_2_2(mux_tmp_687, mux_695_nl, nor_151_cse);
  assign and_381_nl = ((~ operator_3_false_2_operator_3_false_2_and_svs_st_1) | (~
      if_axi_wr_w_PopNB_mioi_bawt) | (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3!=4'b0010))
      & mux_tmp_687;
  assign mux_697_nl = MUX_s_1_2_2(mux_696_nl, and_381_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_698_nl = MUX_s_1_2_2(mux_tmp_687, mux_697_nl, or_dcpl_4);
  assign mux_699_nl = MUX_s_1_2_2(mux_698_nl, mux_tmp_687, or_705_cse);
  assign mux_700_nl = MUX_s_1_2_2(mux_tmp_687, mux_699_nl, or_dcpl_3);
  assign mux_706_nl = MUX_s_1_2_2(mux_tmp_697, mux_tmp_700, regIn_arb_req_sva);
  assign and_393_nl = regIn_arb_req_sva & mux_tmp_700;
  assign nor_157_nl = ~((regIn_PopNB_mioi_idat_mxwt[3:0]!=4'b0001));
  assign mux_707_nl = MUX_s_1_2_2(mux_706_nl, and_393_nl, nor_157_nl);
  assign mux_708_nl = MUX_s_1_2_2(mux_tmp_697, mux_707_nl, nor_151_cse);
  assign nor_302_nl = ~((while_else_4_if_if_regAddr_acc_itm_6_3[0]) | (~ mux_tmp_697));
  assign or_720_nl = (~ operator_3_false_2_operator_3_false_2_and_svs_st_1) | (~
      if_axi_wr_w_PopNB_mioi_bawt) | (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3[3:1]!=3'b000);
  assign mux_703_nl = MUX_s_1_2_2(nor_302_nl, mux_tmp_697, or_720_nl);
  assign mux_709_nl = MUX_s_1_2_2(mux_708_nl, mux_703_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_710_nl = MUX_s_1_2_2(mux_tmp_697, mux_709_nl, or_dcpl_4);
  assign mux_711_nl = MUX_s_1_2_2(mux_710_nl, mux_tmp_697, or_705_cse);
  assign mux_712_nl = MUX_s_1_2_2(mux_tmp_697, mux_711_nl, or_dcpl_3);
  assign and_504_nl = nand_142_cse_1 & (~ mux_725_itm);
  assign and_505_nl = if_axi_rd_r_Push_mioi_bawt & (~ mux_725_itm);
  assign mux_726_nl = MUX_s_1_2_2(and_504_nl, and_505_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign mux_98_nl = MUX_s_1_2_2((~ nand_tmp_10), mux_tmp_86, or_28_cse);
  assign mux_95_nl = MUX_s_1_2_2(nand_tmp_10, (~ nand_tmp_14), while_mux_32_tmp[0]);
  assign or_45_nl = (while_mux_32_tmp[2:1]!=2'b00);
  assign mux_96_nl = MUX_s_1_2_2(mux_95_nl, nand_tmp_10, or_45_nl);
  assign mux_94_nl = MUX_s_1_2_2((~ nand_tmp_10), mux_tmp_86, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_97_nl = MUX_s_1_2_2((~ mux_96_nl), mux_94_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_99_nl = MUX_s_1_2_2(mux_98_nl, mux_97_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_100_nl = MUX_s_1_2_2(mux_99_nl, mux_tmp_86, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_101_nl = MUX_s_1_2_2((~ nand_tmp_10), mux_100_nl, and_309_cse);
  assign mux_89_nl = MUX_s_1_2_2((~ nand_tmp_10), nand_tmp_14, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_90_nl = MUX_s_1_2_2(mux_tmp_86, mux_89_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_91_nl = MUX_s_1_2_2(mux_tmp_87, (~ mux_90_nl), while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign or_74_nl = (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3[3:1]!=3'b100);
  assign mux_92_nl = MUX_s_1_2_2(mux_91_nl, mux_tmp_87, or_74_nl);
  assign mux_93_nl = MUX_s_1_2_2((~ mux_92_nl), mux_tmp_86, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_102_nl = MUX_s_1_2_2(mux_101_nl, mux_93_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nor_nl = ~(mux_102_nl | (~ mux_tmp_724));
  assign mux_731_nl = MUX_s_1_2_2(mux_730_itm, nor_nl, or_dcpl_4);
  assign mux_732_nl = MUX_s_1_2_2(mux_730_itm, mux_731_nl, or_dcpl_2);
  assign mux_733_nl = MUX_s_1_2_2(mux_730_itm, mux_732_nl, or_dcpl_3);
  assign mux_734_nl = MUX_s_1_2_2(mux_733_nl, mux_tmp_724, or_735_cse);
  assign mux_122_nl = MUX_s_1_2_2((~ nand_tmp_15), mux_tmp_112, or_28_cse);
  assign or_27_nl = (while_mux_32_tmp[2:0]!=3'b010);
  assign mux_120_nl = MUX_s_1_2_2(nand_tmp_19, (~ nand_tmp_15), or_27_nl);
  assign mux_119_nl = MUX_s_1_2_2((~ nand_tmp_15), mux_tmp_112, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_121_nl = MUX_s_1_2_2(mux_120_nl, mux_119_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_123_nl = MUX_s_1_2_2(mux_122_nl, mux_121_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_124_nl = MUX_s_1_2_2(mux_123_nl, mux_tmp_112, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_125_nl = MUX_s_1_2_2((~ nand_tmp_15), mux_124_nl, and_309_cse);
  assign mux_115_nl = MUX_s_1_2_2((~ nand_tmp_15), nand_tmp_19, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_116_nl = MUX_s_1_2_2(mux_tmp_112, mux_115_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_113_nl = MUX_s_1_2_2(mux_tmp_112, (~ nand_tmp_15), operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign or_90_nl = (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3!=4'b1010);
  assign mux_117_nl = MUX_s_1_2_2(mux_116_nl, mux_113_nl, or_90_nl);
  assign mux_118_nl = MUX_s_1_2_2(mux_117_nl, mux_tmp_112, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_126_nl = MUX_s_1_2_2(mux_125_nl, mux_118_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nor_387_nl = ~(mux_126_nl | (~ mux_tmp_732));
  assign mux_739_nl = MUX_s_1_2_2(mux_738_itm, nor_387_nl, or_dcpl_4);
  assign mux_740_nl = MUX_s_1_2_2(mux_738_itm, mux_739_nl, or_dcpl_2);
  assign mux_741_nl = MUX_s_1_2_2(mux_738_itm, mux_740_nl, or_dcpl_3);
  assign mux_742_nl = MUX_s_1_2_2(mux_741_nl, mux_tmp_732, or_735_cse);
  assign or_108_nl = (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_6_1) | operator_3_false_1_operator_3_false_1_and_svs_2;
  assign mux_145_nl = MUX_s_1_2_2(mux_tmp_144, mux_tmp_143, or_108_nl);
  assign mux_152_nl = MUX_s_1_2_2(mux_151_cse, mux_145_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_153_nl = MUX_s_1_2_2(or_tmp_103, mux_152_nl, while_stage_v_2);
  assign or_120_nl = (while_mux_32_tmp[1:0]!=2'b10);
  assign mux_154_nl = MUX_s_1_2_2(mux_153_nl, nand_tmp_20, or_120_nl);
  assign mux_155_nl = MUX_s_1_2_2(mux_tmp_149, mux_154_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_150_nl = MUX_s_1_2_2(nand_tmp_20, mux_tmp_149, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_156_nl = MUX_s_1_2_2(mux_155_nl, mux_150_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_157_nl = MUX_s_1_2_2(mux_156_nl, mux_tmp_149, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign nor_133_nl = ~((~((~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_else_4_if_if_for_equal_tmp_6_1) | operator_3_false_1_operator_3_false_1_and_svs_2))
      | mux_5_cse);
  assign mux_138_nl = MUX_s_1_2_2(nor_132_cse, nor_133_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign and_311_nl = while_stage_v_2 & mux_138_nl;
  assign mux_139_nl = MUX_s_1_2_2(nand_tmp_20, and_311_nl, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_140_nl = MUX_s_1_2_2((~ mux_tmp_136), mux_139_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_137_nl = MUX_s_1_2_2((~ mux_tmp_136), nand_tmp_20, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign or_106_nl = (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3!=4'b0110);
  assign mux_141_nl = MUX_s_1_2_2(mux_140_nl, mux_137_nl, or_106_nl);
  assign mux_142_nl = MUX_s_1_2_2(mux_141_nl, (~ mux_tmp_136), operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_158_nl = MUX_s_1_2_2(mux_157_nl, mux_142_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign and_682_nl = mux_158_nl & mux_tmp_740;
  assign mux_747_nl = MUX_s_1_2_2(mux_746_itm, and_682_nl, or_dcpl_4);
  assign mux_748_nl = MUX_s_1_2_2(mux_746_itm, mux_747_nl, or_dcpl_2);
  assign mux_749_nl = MUX_s_1_2_2(mux_746_itm, mux_748_nl, or_dcpl_3);
  assign mux_750_nl = MUX_s_1_2_2(mux_749_nl, mux_tmp_740, or_735_cse);
  assign mux_180_nl = MUX_s_1_2_2((~ nand_tmp_26), mux_tmp_168, or_28_cse);
  assign mux_177_nl = MUX_s_1_2_2(nand_tmp_26, (~ nand_tmp_30), and_312_cse);
  assign mux_178_nl = MUX_s_1_2_2(mux_177_nl, nand_tmp_26, while_mux_32_tmp[2]);
  assign mux_176_nl = MUX_s_1_2_2((~ nand_tmp_26), mux_tmp_168, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_179_nl = MUX_s_1_2_2((~ mux_178_nl), mux_176_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_181_nl = MUX_s_1_2_2(mux_180_nl, mux_179_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_182_nl = MUX_s_1_2_2(mux_181_nl, mux_tmp_168, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_183_nl = MUX_s_1_2_2((~ nand_tmp_26), mux_182_nl, and_309_cse);
  assign mux_171_nl = MUX_s_1_2_2((~ nand_tmp_26), nand_tmp_30, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_172_nl = MUX_s_1_2_2(mux_tmp_168, mux_171_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_173_nl = MUX_s_1_2_2(mux_tmp_169, (~ mux_172_nl), and_314_cse);
  assign or_134_nl = (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3[3:2]!=2'b10);
  assign mux_174_nl = MUX_s_1_2_2(mux_173_nl, mux_tmp_169, or_134_nl);
  assign mux_175_nl = MUX_s_1_2_2((~ mux_174_nl), mux_tmp_168, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_184_nl = MUX_s_1_2_2(mux_183_nl, mux_175_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nor_388_nl = ~(mux_184_nl | (~ mux_tmp_748));
  assign mux_755_nl = MUX_s_1_2_2(mux_754_itm, nor_388_nl, or_dcpl_4);
  assign mux_756_nl = MUX_s_1_2_2(mux_754_itm, mux_755_nl, or_dcpl_2);
  assign mux_757_nl = MUX_s_1_2_2(mux_754_itm, mux_756_nl, or_dcpl_3);
  assign mux_758_nl = MUX_s_1_2_2(mux_757_nl, mux_tmp_748, or_735_cse);
  assign mux_206_nl = MUX_s_1_2_2((~ nand_tmp_31), mux_tmp_194, or_28_cse);
  assign mux_203_nl = MUX_s_1_2_2(nand_tmp_31, (~ nand_tmp_35), and_312_cse);
  assign mux_204_nl = MUX_s_1_2_2(mux_203_nl, nand_tmp_31, while_mux_32_tmp[2]);
  assign mux_202_nl = MUX_s_1_2_2((~ nand_tmp_31), mux_tmp_194, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_205_nl = MUX_s_1_2_2((~ mux_204_nl), mux_202_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_207_nl = MUX_s_1_2_2(mux_206_nl, mux_205_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_208_nl = MUX_s_1_2_2(mux_207_nl, mux_tmp_194, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_209_nl = MUX_s_1_2_2(mux_208_nl, (~ nand_tmp_31), or_26_cse);
  assign mux_197_nl = MUX_s_1_2_2((~ nand_tmp_31), nand_tmp_35, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_198_nl = MUX_s_1_2_2(mux_tmp_194, mux_197_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_199_nl = MUX_s_1_2_2(mux_tmp_195, (~ mux_198_nl), and_314_cse);
  assign or_149_nl = (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3[3:2]!=2'b00);
  assign mux_200_nl = MUX_s_1_2_2(mux_199_nl, mux_tmp_195, or_149_nl);
  assign mux_201_nl = MUX_s_1_2_2((~ mux_200_nl), mux_tmp_194, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_210_nl = MUX_s_1_2_2(mux_209_nl, mux_201_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nor_389_nl = ~(mux_210_nl | (~ mux_tmp_756));
  assign mux_763_nl = MUX_s_1_2_2(mux_762_itm, nor_389_nl, or_dcpl_4);
  assign mux_764_nl = MUX_s_1_2_2(mux_762_itm, mux_763_nl, or_dcpl_2);
  assign mux_765_nl = MUX_s_1_2_2(mux_762_itm, mux_764_nl, or_dcpl_3);
  assign mux_766_nl = MUX_s_1_2_2(mux_765_nl, mux_tmp_756, or_735_cse);
  assign nand_195_nl = ~(while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1
      & while_else_4_if_if_for_equal_tmp_7_1);
  assign mux_230_nl = MUX_s_1_2_2(mux_tmp_144, mux_tmp_143, nand_195_nl);
  assign mux_237_nl = MUX_s_1_2_2(mux_151_cse, mux_230_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_239_nl = MUX_s_1_2_2(nand_tmp_36, mux_237_nl, and_312_cse);
  assign mux_240_nl = MUX_s_1_2_2(mux_tmp_234, mux_239_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_235_nl = MUX_s_1_2_2(nand_tmp_36, mux_tmp_234, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_241_nl = MUX_s_1_2_2(mux_240_nl, mux_235_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_242_nl = MUX_s_1_2_2(mux_241_nl, mux_tmp_234, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign nor_135_nl = ~(and_499_cse | mux_5_cse);
  assign mux_222_nl = MUX_s_1_2_2(nor_132_cse, nor_135_nl, operator_3_false_2_operator_3_false_2_and_svs_2);
  assign mux_223_nl = MUX_s_1_2_2(nand_tmp_36, mux_222_nl, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_224_nl = MUX_s_1_2_2((~ mux_tmp_220), mux_223_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign and_318_nl = (while_else_4_if_if_regAddr_acc_itm_6_3[2:0]==3'b111);
  assign mux_225_nl = MUX_s_1_2_2(mux_tmp_221, mux_224_nl, and_318_nl);
  assign or_165_nl = (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3[3]);
  assign mux_226_nl = MUX_s_1_2_2(mux_225_nl, mux_tmp_221, or_165_nl);
  assign mux_227_nl = MUX_s_1_2_2(mux_226_nl, (~ mux_tmp_220), operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_243_nl = MUX_s_1_2_2(mux_242_nl, mux_227_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign and_683_nl = mux_243_nl & mux_tmp_764;
  assign mux_771_nl = MUX_s_1_2_2(mux_770_itm, and_683_nl, or_dcpl_4);
  assign mux_772_nl = MUX_s_1_2_2(mux_770_itm, mux_771_nl, or_dcpl_2);
  assign mux_773_nl = MUX_s_1_2_2(mux_770_itm, mux_772_nl, or_dcpl_3);
  assign mux_774_nl = MUX_s_1_2_2(mux_773_nl, mux_tmp_764, or_735_cse);
  assign mux_263_nl = MUX_s_1_2_2((~ nand_tmp_42), mux_tmp_253, or_28_cse);
  assign or_194_nl = (while_mux_32_tmp[2:0]!=3'b100);
  assign mux_261_nl = MUX_s_1_2_2(nand_tmp_46, (~ nand_tmp_42), or_194_nl);
  assign mux_260_nl = MUX_s_1_2_2((~ nand_tmp_42), mux_tmp_253, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_262_nl = MUX_s_1_2_2(mux_261_nl, mux_260_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_264_nl = MUX_s_1_2_2(mux_263_nl, mux_262_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_265_nl = MUX_s_1_2_2(mux_264_nl, mux_tmp_253, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_266_nl = MUX_s_1_2_2((~ nand_tmp_42), mux_265_nl, and_309_cse);
  assign mux_256_nl = MUX_s_1_2_2((~ nand_tmp_42), nand_tmp_46, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_257_nl = MUX_s_1_2_2(mux_tmp_253, mux_256_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_254_nl = MUX_s_1_2_2(mux_tmp_253, (~ nand_tmp_42), operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign or_192_nl = (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3!=4'b1100);
  assign mux_258_nl = MUX_s_1_2_2(mux_257_nl, mux_254_nl, or_192_nl);
  assign mux_259_nl = MUX_s_1_2_2(mux_258_nl, mux_tmp_253, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_267_nl = MUX_s_1_2_2(mux_266_nl, mux_259_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nor_390_nl = ~(mux_267_nl | (~ mux_tmp_772));
  assign mux_779_nl = MUX_s_1_2_2(mux_778_itm, nor_390_nl, or_dcpl_4);
  assign mux_780_nl = MUX_s_1_2_2(mux_778_itm, mux_779_nl, or_dcpl_2);
  assign mux_781_nl = MUX_s_1_2_2(mux_778_itm, mux_780_nl, or_dcpl_3);
  assign mux_782_nl = MUX_s_1_2_2(mux_781_nl, mux_tmp_772, or_735_cse);
  assign mux_289_nl = MUX_s_1_2_2((~ nand_tmp_47), mux_tmp_277, or_28_cse);
  assign mux_286_nl = MUX_s_1_2_2(nand_tmp_47, (~ nand_tmp_51), while_mux_32_tmp[0]);
  assign mux_287_nl = MUX_s_1_2_2(mux_286_nl, nand_tmp_47, or_210_cse);
  assign mux_285_nl = MUX_s_1_2_2((~ nand_tmp_47), mux_tmp_277, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_288_nl = MUX_s_1_2_2((~ mux_287_nl), mux_285_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_290_nl = MUX_s_1_2_2(mux_289_nl, mux_288_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_291_nl = MUX_s_1_2_2(mux_290_nl, mux_tmp_277, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_292_nl = MUX_s_1_2_2((~ nand_tmp_47), mux_291_nl, and_309_cse);
  assign mux_280_nl = MUX_s_1_2_2((~ nand_tmp_47), nand_tmp_51, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_281_nl = MUX_s_1_2_2(mux_tmp_277, mux_280_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_282_nl = MUX_s_1_2_2(mux_tmp_278, (~ mux_281_nl), while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign nand_143_nl = ~(if_axi_wr_w_PopNB_mioi_ivld_mxwt & (while_else_4_if_if_regAddr_acc_itm_6_3[3:1]==3'b110));
  assign mux_283_nl = MUX_s_1_2_2(mux_282_nl, mux_tmp_278, nand_143_nl);
  assign mux_284_nl = MUX_s_1_2_2((~ mux_283_nl), mux_tmp_277, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_293_nl = MUX_s_1_2_2(mux_292_nl, mux_284_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nor_391_nl = ~(mux_293_nl | (~ mux_tmp_780));
  assign mux_787_nl = MUX_s_1_2_2(mux_786_itm, nor_391_nl, or_dcpl_4);
  assign mux_788_nl = MUX_s_1_2_2(mux_786_itm, mux_787_nl, or_dcpl_2);
  assign mux_789_nl = MUX_s_1_2_2(mux_786_itm, mux_788_nl, or_dcpl_3);
  assign mux_790_nl = MUX_s_1_2_2(mux_789_nl, mux_tmp_780, or_735_cse);
  assign mux_315_nl = MUX_s_1_2_2((~ nand_tmp_52), mux_tmp_303, or_28_cse);
  assign mux_312_nl = MUX_s_1_2_2(nand_tmp_52, (~ nand_tmp_56), while_mux_32_tmp[0]);
  assign mux_313_nl = MUX_s_1_2_2(mux_312_nl, nand_tmp_52, or_210_cse);
  assign mux_311_nl = MUX_s_1_2_2((~ nand_tmp_52), mux_tmp_303, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_314_nl = MUX_s_1_2_2((~ mux_313_nl), mux_311_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_316_nl = MUX_s_1_2_2(mux_315_nl, mux_314_nl, operator_3_false_3_operator_3_false_3_and_svs_st_1);
  assign mux_317_nl = MUX_s_1_2_2(mux_316_nl, mux_tmp_303, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_318_nl = MUX_s_1_2_2(mux_317_nl, (~ nand_tmp_52), or_26_cse);
  assign mux_306_nl = MUX_s_1_2_2((~ nand_tmp_52), nand_tmp_56, if_axi_wr_w_PopNB_mioi_bawt);
  assign mux_307_nl = MUX_s_1_2_2(mux_tmp_303, mux_306_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_308_nl = MUX_s_1_2_2(mux_tmp_304, (~ mux_307_nl), while_else_4_if_if_regAddr_acc_itm_6_3[0]);
  assign or_224_nl = (~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) | (while_else_4_if_if_regAddr_acc_itm_6_3[3:1]!=3'b010);
  assign mux_309_nl = MUX_s_1_2_2(mux_308_nl, mux_tmp_304, or_224_nl);
  assign mux_310_nl = MUX_s_1_2_2((~ mux_309_nl), mux_tmp_303, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_319_nl = MUX_s_1_2_2(mux_318_nl, mux_310_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign nor_392_nl = ~(mux_319_nl | (~ mux_tmp_788));
  assign mux_795_nl = MUX_s_1_2_2(mux_794_itm, nor_392_nl, or_dcpl_4);
  assign mux_796_nl = MUX_s_1_2_2(mux_794_itm, mux_795_nl, or_dcpl_2);
  assign mux_797_nl = MUX_s_1_2_2(mux_794_itm, mux_796_nl, or_dcpl_3);
  assign mux_798_nl = MUX_s_1_2_2(mux_797_nl, mux_tmp_788, or_735_cse);
  assign while_else_4_mux_20_nl = MUX_s_1_2_2(while_else_4_else_while_else_4_else_and_itm,
      while_while_or_2_tmp, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign while_else_4_if_mux_17_nl = MUX_s_1_2_2(while_while_or_1_tmp, while_else_4_if_if_while_else_4_if_if_and_1_itm,
      if_axi_wr_w_PopNB_mioi_ivld_mxwt);
  assign while_else_4_mux_22_nl = MUX_s_1_2_2(while_while_or_1_tmp, while_else_4_if_mux_17_nl,
      operator_3_false_2_operator_3_false_2_and_svs_1);
  assign while_if_4_while_if_4_or_1_nl = arb_needs_update_sva | operator_8_false_operator_8_false_nor_mdf_sva_mx1;
  assign while_else_4_else_while_else_4_else_or_nl = arb_needs_update_sva | operator_3_false_3_operator_3_false_3_and_svs_1;
  assign while_else_4_if_if_while_else_4_if_if_or_nl = arb_needs_update_sva | (if_axi_wr_w_PopNB_mioi_idat_mxwt[64]);
  assign while_if_4_nand_nl = ~((~((~ if_axi_wr_w_PopNB_mioi_ivld_mxwt) & while_and_110_cse))
      & while_stage_v_1);
  assign while_if_4_mux1h_3_nl = MUX1HOT_s_1_4_2(while_if_4_while_if_4_or_1_nl, while_else_4_else_while_else_4_else_or_nl,
      arb_needs_update_sva, while_else_4_if_if_while_else_4_if_if_or_nl, {and_dcpl_77
      , while_if_4_and_1_cse , while_if_4_nand_nl , while_if_4_and_4_cse});
  assign nl_while_if_4_else_2_acc_nl = axiRdLen_sva_dfm_1_mx0 + 8'b11111111;
  assign while_if_4_else_2_acc_nl = nl_while_if_4_else_2_acc_nl[7:0];
  assign nor_128_nl = ~((~ if_axi_wr_w_PopNB_mioi_bawt) | (if_axi_wr_w_PopNB_mioi_idat_mxwt[64])
      | (~(if_axi_wr_w_PopNB_mioi_ivld_mxwt & or_dcpl_25)));
  assign mux_501_nl = MUX_s_1_2_2(or_dcpl_25, nor_128_nl, nor_tmp_28);
  assign nand_172_nl = ~(or_28_cse & or_dcpl_25);
  assign or_486_nl = while_if_4_aelse_acc_itm_16_1 | while_if_4_acc_1_itm_16_1 |
      and_dcpl_35;
  assign mux_506_nl = MUX_s_1_2_2(nand_172_nl, or_486_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign and_167_nl = or_tmp_435 & or_dcpl_25;
  assign mux_547_nl = MUX_s_1_2_2((~ or_tmp_287), or_dcpl_25, nor_tmp_30);
  assign mux_546_nl = MUX_s_1_2_2((~ or_tmp_287), or_dcpl_25, or_tmp_439);
  assign mux_548_nl = MUX_s_1_2_2(mux_547_nl, mux_546_nl, arb_next_1_1_sva);
  assign mux_549_nl = MUX_s_1_2_2(and_167_nl, mux_548_nl, arb_needs_update_sva);
  assign mux_550_nl = MUX_s_1_2_2(mux_549_nl, mux_tmp_545, while_stage_v_1);
  assign while_or_25_nl = and_dcpl_79 | while_and_104_cse;
  assign while_or_26_nl = and_dcpl_79 | while_and_103_cse | ((~ if_axi_wr_w_PopNB_mioi_ivld_mxwt)
      & while_and_104_cse);
  assign while_and_108_nl = if_axi_wr_w_PopNB_mioi_ivld_mxwt & while_and_104_cse;
  assign nand_144_nl = ~((operator_3_false_1_operator_3_false_1_and_svs_2 | (~ while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ operator_3_false_2_operator_3_false_2_and_svs_2) | while_else_4_if_if_while_else_4_if_if_nand_tmp_1)
      & operator_3_false_2_operator_3_false_2_and_svs_st_2 & while_else_4_if_Connections_InBlocking_axi_axi4_axi_cfg_standard_WritePayload_Connections_SYN_PORT_PopNB_return_sva_st_1
      & while_else_4_if_if_slc_if_axi_wr_w_PopNB_mio_mrgout_dat_64_itm_1 & (~ if_axi_wr_b_Push_mioi_bawt));
  assign mux_331_nl = MUX_s_1_2_2(nand_144_nl, if_axi_rd_r_Push_mioi_bawt, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign and_323_nl = while_stage_v_2 & (~ mux_331_nl);
  assign mux_332_nl = MUX_s_1_2_2(or_tmp_228, and_323_nl, or_dcpl_3);
  assign mux_333_nl = MUX_s_1_2_2(or_tmp_228, mux_332_nl, or_dcpl_2);
  assign and_322_nl = operator_3_false_2_operator_3_false_2_and_svs_st_1 & (if_axi_wr_w_PopNB_mioi_idat_mxwt[72:65]==8'b11111111)
      & if_axi_wr_w_PopNB_mioi_ivld_mxwt & if_axi_wr_w_PopNB_mioi_bawt;
  assign mux_334_nl = MUX_s_1_2_2(or_tmp_228, mux_333_nl, and_322_nl);
  assign or_248_nl = (~ or_dcpl_4) | (~ while_stage_v_1) | operator_3_false_1_operator_3_false_1_and_svs_1
      | (~ operator_3_false_2_operator_3_false_2_and_svs_1) | operator_3_false_1_operator_3_false_1_and_svs_st_1;
  assign mux_335_nl = MUX_s_1_2_2(mux_334_nl, or_tmp_228, or_248_nl);
  assign nand_208_nl = ~(nand_142_cse_1 & or_tmp_762);
  assign nand_209_nl = ~(if_axi_rd_r_Push_mioi_bawt & or_tmp_762);
  assign mux_834_nl = MUX_s_1_2_2(nand_208_nl, nand_209_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nand_212_nl = ~(nand_142_cse_1 & or_tmp_778);
  assign nand_213_nl = ~(if_axi_rd_r_Push_mioi_bawt & or_tmp_778);
  assign mux_850_nl = MUX_s_1_2_2(nand_212_nl, nand_213_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign nand_216_nl = ~(nand_142_cse_1 & or_tmp_794);
  assign nand_217_nl = ~(if_axi_rd_r_Push_mioi_bawt & or_tmp_794);
  assign mux_866_nl = MUX_s_1_2_2(nand_216_nl, nand_217_nl, operator_3_false_1_operator_3_false_1_and_svs_st_2);
  assign and_189_nl = or_dcpl_64 & (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[69]));
  assign and_191_nl = or_dcpl_64 & (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[68]));
  assign and_193_nl = or_dcpl_64 & (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[67]));
  assign and_195_nl = or_dcpl_64 & (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[66]));
  assign and_197_nl = or_dcpl_64 & (~ (if_axi_wr_w_PopNB_mioi_idat_mxwt[65]));
  assign nand_109_nl = ~(select_mask_2_1_sva_1 & (~(arb_next_1_1_sva & write_arb_req_sva))
      & nand_tmp_98);
  assign or_602_nl = select_mask_2_1_sva_1 | nor_tmp_30 | (~ nand_tmp_98);
  assign mux_673_nl = MUX_s_1_2_2(nand_109_nl, or_602_nl, select_mask_2_1_sva_0);
  assign or_600_nl = (regIn_arb_req_sva & write_arb_req_sva) | read_arb_req_sva |
      (~ nand_tmp_98);
  assign mux_670_nl = MUX_s_1_2_2(or_tmp_510, or_tmp_529, regIn_arb_req_sva);
  assign mux_671_nl = MUX_s_1_2_2(or_600_nl, mux_670_nl, arb_next_1_2_sva);
  assign mux_668_nl = MUX_s_1_2_2(or_tmp_510, (~ nand_tmp_98), write_arb_req_sva);
  assign mux_669_nl = MUX_s_1_2_2(mux_668_nl, or_tmp_529, nor_tmp_30);
  assign mux_672_nl = MUX_s_1_2_2(mux_671_nl, mux_669_nl, arb_next_1_1_sva);
  assign mux_674_nl = MUX_s_1_2_2(mux_673_nl, mux_672_nl, arb_needs_update_sva);
  assign mux_665_nl = MUX_s_1_2_2(not_tmp_373, mux_tmp_656, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign mux_657_nl = MUX_s_1_2_2(nand_tmp_103, (~ and_tmp_75), regIn_PopNB_mioi_ivld_mxwt);
  assign mux_658_nl = MUX_s_1_2_2(mux_657_nl, nand_tmp_102, while_asn_34_itm_1);
  assign mux_659_nl = MUX_s_1_2_2((~ mux_658_nl), and_tmp_76, regIn_arb_req_sva);
  assign mux_660_nl = MUX_s_1_2_2(not_tmp_372, mux_659_nl, arb_next_1_2_sva);
  assign mux_662_nl = MUX_s_1_2_2((~ mux_tmp_633), mux_660_nl, and_352_cse);
  assign mux_663_nl = MUX_s_1_2_2(mux_tmp_653, mux_662_nl, operator_3_false_2_operator_3_false_2_and_svs_1);
  assign mux_664_nl = MUX_s_1_2_2(mux_663_nl, (~ mux_tmp_656), operator_3_false_1_operator_3_false_1_and_svs_1);
  assign nand_108_nl = ~(if_axi_wr_w_PopNB_mioi_bawt & mux_664_nl);
  assign mux_666_nl = MUX_s_1_2_2(mux_665_nl, nand_108_nl, operator_3_false_2_operator_3_false_2_and_svs_st_1);
  assign mux_643_nl = MUX_s_1_2_2(mux_tmp_642, mux_tmp_633, or_310_cse);
  assign mux_655_nl = MUX_s_1_2_2(not_tmp_373, mux_643_nl, operator_3_false_1_operator_3_false_1_and_svs_1);
  assign mux_667_nl = MUX_s_1_2_2(mux_666_nl, mux_655_nl, operator_3_false_1_operator_3_false_1_and_svs_st_1);
  assign mux_675_nl = MUX_s_1_2_2(mux_674_nl, mux_667_nl, while_stage_v_1);
  assign mux_676_nl = MUX_s_1_2_2(or_dcpl_25, and_dcpl_26, while_stage_v_1);
  assign while_else_4_if_if_aelse_mux_2_nl = MUX_v_16_2_2(operator_33_true_return_15_0_sva,
      baseAddr, fsm_output[0]);
  assign while_else_4_if_if_aelse_or_1_nl = (fsm_output!=2'b01);
  assign while_else_4_if_if_aelse_mux_3_nl = MUX_v_13_2_2((~ axiWrAddr_15_3_sva_dfm_1_mx0),
      13'b0000000001101, fsm_output[0]);
  assign while_else_4_if_if_aelse_not_1_nl = ~ (fsm_output[0]);
  assign while_else_4_if_if_aelse_while_else_4_if_if_aelse_while_else_4_if_if_aelse_nand_1_nl
      = ~(MUX_v_3_2_2(3'b000, axiWrAddr_2_0_sva_dfm_1_mx1, while_else_4_if_if_aelse_not_1_nl));
  assign nl_acc_nl = ({(~ (fsm_output[0])) , while_else_4_if_if_aelse_mux_2_nl ,
      while_else_4_if_if_aelse_or_1_nl}) + conv_u2u_17_18({while_else_4_if_if_aelse_mux_3_nl
      , while_else_4_if_if_aelse_while_else_4_if_if_aelse_while_else_4_if_if_aelse_nand_1_nl
      , 1'b1});
  assign acc_nl = nl_acc_nl[17:0];
  assign z_out = readslicef_18_17_1(acc_nl);
  assign and_684_nl = (~ operator_3_false_1_operator_3_false_1_and_svs_1) & (fsm_output[1]);
  assign operator_16_false_mux_1_nl = MUX_v_13_2_2(axiRdAddr_15_3_sva_dfm_1_mx0,
      axiWrAddr_15_3_sva_dfm_1_mx0, and_684_nl);
  assign nl_z_out_1 = operator_16_false_mux_1_nl + 13'b0000000000001;
  assign z_out_1 = nl_z_out_1[12:0];

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | (input_1 & {64{sel[1]}});
    result = result | (input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_14_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [63:0] input_2;
    input [63:0] input_3;
    input [63:0] input_4;
    input [63:0] input_5;
    input [63:0] input_6;
    input [63:0] input_7;
    input [63:0] input_8;
    input [63:0] input_9;
    input [63:0] input_10;
    input [63:0] input_11;
    input [63:0] input_12;
    input [63:0] input_13;
    input [3:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      default : begin
        result = input_13;
      end
    endcase
    MUX_v_64_14_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction


  function automatic [3:0] readslicef_7_4_3;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_7_4_3 = tmp[3:0];
  end
  endfunction


  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_u2u_17_18 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AxiSlaveToReg2_axi_cfg_standard_14_16
// ------------------------------------------------------------------


module AxiSlaveToReg2_axi_cfg_standard_14_16 (
  clk, reset_bar, if_axi_rd_ar_val, if_axi_rd_ar_rdy, if_axi_rd_ar_msg, if_axi_rd_r_val,
      if_axi_rd_r_rdy, if_axi_rd_r_msg, if_axi_wr_aw_val, if_axi_wr_aw_rdy, if_axi_wr_aw_msg,
      if_axi_wr_w_val, if_axi_wr_w_rdy, if_axi_wr_w_msg, if_axi_wr_b_val, if_axi_wr_b_rdy,
      if_axi_wr_b_msg, baseAddr, regOut_0, regOut_1, regOut_2, regOut_3, regOut_4,
      regOut_5, regOut_6, regOut_7, regOut_8, regOut_9, regOut_10, regOut_11, regOut_12,
      regOut_13, regIn_val, regIn_rdy, regIn_msg
);
  input clk;
  input reset_bar;
  input if_axi_rd_ar_val;
  output if_axi_rd_ar_rdy;
  input [43:0] if_axi_rd_ar_msg;
  output if_axi_rd_r_val;
  input if_axi_rd_r_rdy;
  output [70:0] if_axi_rd_r_msg;
  input if_axi_wr_aw_val;
  output if_axi_wr_aw_rdy;
  input [43:0] if_axi_wr_aw_msg;
  input if_axi_wr_w_val;
  output if_axi_wr_w_rdy;
  input [72:0] if_axi_wr_w_msg;
  output if_axi_wr_b_val;
  input if_axi_wr_b_rdy;
  output [5:0] if_axi_wr_b_msg;
  input [15:0] baseAddr;
  output [63:0] regOut_0;
  output [63:0] regOut_1;
  output [63:0] regOut_2;
  output [63:0] regOut_3;
  output [63:0] regOut_4;
  output [63:0] regOut_5;
  output [63:0] regOut_6;
  output [63:0] regOut_7;
  output [63:0] regOut_8;
  output [63:0] regOut_9;
  output [63:0] regOut_10;
  output [63:0] regOut_11;
  output [63:0] regOut_12;
  output [63:0] regOut_13;
  input regIn_val;
  output regIn_rdy;
  input [70:0] regIn_msg;



  // Interconnect Declarations for Component Instantiations 
  AxiSlaveToReg2_axi_cfg_standard_14_16_run AxiSlaveToReg2_axi_cfg_standard_14_16_run_inst
      (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_rd_ar_val(if_axi_rd_ar_val),
      .if_axi_rd_ar_rdy(if_axi_rd_ar_rdy),
      .if_axi_rd_ar_msg(if_axi_rd_ar_msg),
      .if_axi_rd_r_val(if_axi_rd_r_val),
      .if_axi_rd_r_rdy(if_axi_rd_r_rdy),
      .if_axi_rd_r_msg(if_axi_rd_r_msg),
      .if_axi_wr_aw_val(if_axi_wr_aw_val),
      .if_axi_wr_aw_rdy(if_axi_wr_aw_rdy),
      .if_axi_wr_aw_msg(if_axi_wr_aw_msg),
      .if_axi_wr_w_val(if_axi_wr_w_val),
      .if_axi_wr_w_rdy(if_axi_wr_w_rdy),
      .if_axi_wr_w_msg(if_axi_wr_w_msg),
      .if_axi_wr_b_val(if_axi_wr_b_val),
      .if_axi_wr_b_rdy(if_axi_wr_b_rdy),
      .if_axi_wr_b_msg(if_axi_wr_b_msg),
      .baseAddr(baseAddr),
      .regOut_0(regOut_0),
      .regOut_1(regOut_1),
      .regOut_2(regOut_2),
      .regOut_3(regOut_3),
      .regOut_4(regOut_4),
      .regOut_5(regOut_5),
      .regOut_6(regOut_6),
      .regOut_7(regOut_7),
      .regOut_8(regOut_8),
      .regOut_9(regOut_9),
      .regOut_10(regOut_10),
      .regOut_11(regOut_11),
      .regOut_12(regOut_12),
      .regOut_13(regOut_13),
      .regIn_val(regIn_val),
      .regIn_rdy(regIn_rdy),
      .regIn_msg(regIn_msg)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Accelerator_rtl
// ------------------------------------------------------------------


module Accelerator_rtl (
  clk, reset_bar, axi_read_ar_val, axi_read_ar_rdy, axi_read_ar_msg, axi_read_r_val,
      axi_read_r_rdy, axi_read_r_msg, axi_write_aw_val, axi_write_aw_rdy, axi_write_aw_msg,
      axi_write_w_val, axi_write_w_rdy, axi_write_w_msg, axi_write_b_val, axi_write_b_rdy,
      axi_write_b_msg
);
  input clk;
  input reset_bar;
  input axi_read_ar_val;
  output axi_read_ar_rdy;
  input [43:0] axi_read_ar_msg;
  output axi_read_r_val;
  input axi_read_r_rdy;
  output [70:0] axi_read_r_msg;
  input axi_write_aw_val;
  output axi_write_aw_rdy;
  input [43:0] axi_write_aw_msg;
  input axi_write_w_val;
  output axi_write_w_rdy;
  input [72:0] axi_write_w_msg;
  output axi_write_b_val;
  input axi_write_b_rdy;
  output [5:0] axi_write_b_msg;


  // Interconnect Declarations
  wire [63:0] regOut_chan_0;
  wire [63:0] regOut_chan_1;
  wire [63:0] regOut_chan_2;
  wire [63:0] regOut_chan_3;
  wire [63:0] regOut_chan_4;
  wire [63:0] regOut_chan_5;
  wire [63:0] regOut_chan_6;
  wire [63:0] regOut_chan_7;
  wire [63:0] regOut_chan_8;
  wire [63:0] regOut_chan_9;
  wire [63:0] regOut_chan_10;
  wire [63:0] regOut_chan_11;
  wire [63:0] regOut_chan_12;
  wire [63:0] regOut_chan_13;
  wire regIn_chan_val;
  wire regIn_chan_rdy;
  wire [70:0] regIn_chan_msg;


  // Interconnect Declarations for Component Instantiations 
  AxiSlaveToReg2_axi_cfg_standard_14_16 slave (
      .clk(clk),
      .reset_bar(reset_bar),
      .if_axi_rd_ar_val(axi_read_ar_val),
      .if_axi_rd_ar_rdy(axi_read_ar_rdy),
      .if_axi_rd_ar_msg(axi_read_ar_msg),
      .if_axi_rd_r_val(axi_read_r_val),
      .if_axi_rd_r_rdy(axi_read_r_rdy),
      .if_axi_rd_r_msg(axi_read_r_msg),
      .if_axi_wr_aw_val(axi_write_aw_val),
      .if_axi_wr_aw_rdy(axi_write_aw_rdy),
      .if_axi_wr_aw_msg(axi_write_aw_msg),
      .if_axi_wr_w_val(axi_write_w_val),
      .if_axi_wr_w_rdy(axi_write_w_rdy),
      .if_axi_wr_w_msg(axi_write_w_msg),
      .if_axi_wr_b_val(axi_write_b_val),
      .if_axi_wr_b_rdy(axi_write_b_rdy),
      .if_axi_wr_b_msg(axi_write_b_msg),
      .baseAddr(16'b0000000000000000),
      .regOut_0(regOut_chan_0),
      .regOut_1(regOut_chan_1),
      .regOut_2(regOut_chan_2),
      .regOut_3(regOut_chan_3),
      .regOut_4(regOut_chan_4),
      .regOut_5(regOut_chan_5),
      .regOut_6(regOut_chan_6),
      .regOut_7(regOut_chan_7),
      .regOut_8(regOut_chan_8),
      .regOut_9(regOut_chan_9),
      .regOut_10(regOut_chan_10),
      .regOut_11(regOut_chan_11),
      .regOut_12(regOut_chan_12),
      .regOut_13(regOut_chan_13),
      .regIn_val(regIn_chan_val),
      .regIn_rdy(regIn_chan_rdy),
      .regIn_msg(regIn_chan_msg)
    );
  Accelerator_run Accelerator_inst (
      .clk(clk),
      .reset_bar(reset_bar),
      .regOut_chan_0(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .regOut_chan_1(regOut_chan_1),
      .regOut_chan_2(regOut_chan_2),
      .regOut_chan_3(regOut_chan_3),
      .regOut_chan_4(regOut_chan_4),
      .regOut_chan_5(regOut_chan_5),
      .regOut_chan_6(regOut_chan_6),
      .regOut_chan_7(regOut_chan_7),
      .regOut_chan_8(regOut_chan_8),
      .regOut_chan_9(regOut_chan_9),
      .regIn_chan_val(regIn_chan_val),
      .regIn_chan_rdy(regIn_chan_rdy),
      .regIn_chan_msg(regIn_chan_msg)
    );
endmodule



